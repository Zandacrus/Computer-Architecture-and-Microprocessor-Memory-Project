

package MATRIX_MULTIPLY_32_PKG;
	
	import MATRIX_MULTIPLY_32_PKG_7::DATA7;
	
	parameter MM32_DATA_SIZE = 67235, SIZE_LIMIT = 8500;
	
	int DATA0 [MM32_DATA_SIZE-(7*SIZE_LIMIT)-1:0] = {'h10b4c, 'h107ac, 'h10944, 'h107bc, 'h107cc, 'h10945, 'h107dc, 'h107ec, 'h10946, 'h107fc, 'h1080c, 'h10947, 'h1081c, 'h103bc, 'h1082c, 'h10948, 'h1083c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084c, 'h10949, 'h10b4c, 'h1085c, 'h1086c, 'h1094a, 'h1087c, 'h1088c, 'h1094b, 'h1089c, 'h108ac, 'h1094c, 'h108bc, 'h108cc, 'h1094d, 'h103bc, 'h108dc, 'h106ec, 'h1094e, 'h10b5c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fc, 'h1070c, 'h1094f, 'h1071c, 'h1072c, 'h10950, 'h1073c, 'h1074c, 'h10951, 'h1075c, 'h1076c, 'h10952, 'h1077c, 'h103bc, 'h1078c, 'h10953, 'h1079c, 'h10b5c, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ac, 'h10954, 'h107bc, 'h107cc, 'h10955, 'h107dc, 'h107ec, 'h10956, 'h107fc, 'h1080c, 'h10957, 'h1081c, 'h1082c, 'h10958, 'h103bc, 'h1083c, 'h1084c, 'h10959, 'h10b5c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085c, 'h1086c, 'h1095a, 'h1087c, 'h1088c, 'h1095b, 'h1089c, 'h108ac, 'h1095c, 'h108bc, 'h108cc, 'h1095d, 'h108dc, 'h103bc, 'h106ec, 'h1095e, 'h10b6c, 'h106fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h1095f, 'h1071c, 'h1072c, 'h10960, 'h1073c, 'h1074c, 'h10961, 'h1075c, 'h1076c, 'h10962, 'h1077c, 'h1078c, 'h10963, 'h103bc, 'h1079c, 'h10b6c, 'h107ac, 'h10964, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bc, 'h107cc, 'h10965, 'h107dc, 'h107ec, 'h10966, 'h107fc, 'h1080c, 'h10967, 'h1081c, 'h1082c, 'h10968, 'h1083c, 'h103bc, 'h1084c, 'h10969, 'h10b6c, 'h1085c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086c, 'h1096a, 'h1087c, 'h1088c, 'h1096b, 'h1089c, 'h108ac, 'h1096c, 'h108bc, 'h108cc, 'h1096d, 'h108dc, 'h106ec, 'h1096e, 'h10b7c, 'h103bc, 'h106fc, 'h1070c, 'h1096f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071c, 'h1072c, 'h10970, 'h1073c, 'h1074c, 'h10971, 'h1075c, 'h1076c, 'h10972, 'h1077c, 'h1078c, 'h10973, 'h1079c, 'h10b7c, 'h103bc, 'h107ac, 'h10974, 'h107bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cc, 'h10975, 'h107dc, 'h107ec, 'h10976, 'h107fc, 'h1080c, 'h10977, 'h1081c, 'h1082c, 'h10978, 'h1083c, 'h1084c, 'h10979, 'h10b7c, 'h103bc, 'h1085c, 'h1086c, 'h1097a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087c, 'h1088c, 'h1097b, 'h1089c, 'h108ac, 'h1097c, 'h108bc, 'h108cc, 'h1097d, 'h108dc, 'h106ec, 'h1097e, 'h10b8c, 'h106fc, 'h103bc, 'h1070c, 'h1097f, 'h1071c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072c, 'h10980, 'h1073c, 'h1074c, 'h10981, 'h1075c, 'h1076c, 'h10982, 'h1077c, 'h1078c, 'h10983, 'h1079c, 'h10b8c, 'h107ac, 'h10984, 'h103bc, 'h107bc, 'h107cc, 'h10985, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dc, 'h107ec, 'h10986, 'h107fc, 'h1080c, 'h10987, 'h1081c, 'h1082c, 'h10988, 'h1083c, 'h1084c, 'h10989, 'h10b8c, 'h1085c, 'h103bc, 'h1086c, 'h1098a, 'h1087c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088c, 'h1098b, 'h1089c, 'h108ac, 'h1098c, 'h108bc, 'h108cc, 'h1098d, 'h108dc, 'h106ec, 'h1098e, 'h10b9c, 'h106fc, 'h1070c, 'h1098f, 'h103bc, 'h1071c, 'h1072c, 'h10990, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h1074c, 'h10991, 'h1075c, 'h1076c, 'h10992, 'h1077c, 'h1078c, 'h10993, 'h1079c, 'h10b9c, 'h107ac, 'h10994, 'h107bc, 'h103bc, 'h107cc, 'h10995, 'h107dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ec, 'h10996, 'h107fc, 'h1080c, 'h10997, 'h1081c, 'h1082c, 'h10998, 'h1083c, 'h1084c, 'h10999, 'h10b9c, 'h1085c, 'h1086c, 'h1099a, 'h103bc, 'h1087c, 'h1088c, 'h1099b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089c, 'h108ac, 'h1099c, 'h108bc, 'h108cc, 'h1099d, 'h108dc, 'h106ec, 'h1099e, 'h10bac, 'h106fc, 'h1070c, 'h1099f, 'h1071c, 'h103bc, 'h1072c, 'h109a0, 'h1073c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074c, 'h109a1, 'h1075c, 'h1076c, 'h109a2, 'h1077c, 'h1078c, 'h109a3, 'h1079c, 'h10bac, 'h107ac, 'h109a4, 'h107bc, 'h107cc, 'h109a5, 'h103bc, 'h107dc, 'h107ec, 'h109a6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fc, 'h1080c, 'h109a7, 'h1081c, 'h1082c, 'h109a8, 'h1083c, 'h1084c, 'h109a9, 'h10bac, 'h1085c, 'h1086c, 'h109aa, 'h1087c, 'h103bc, 'h1088c, 'h109ab, 'h1089c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ac, 'h109ac, 'h108bc, 'h108cc, 'h109ad, 'h108dc, 'h106ec, 'h109ae, 'h10bbc, 'h106fc, 'h1070c, 'h109af, 'h1071c, 'h1072c, 'h109b0, 'h103bc, 'h1073c, 'h1074c, 'h109b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075c, 'h1076c, 'h109b2, 'h1077c, 'h1078c, 'h109b3, 'h1079c, 'h10bbc, 'h107ac, 'h109b4, 'h107bc, 'h107cc, 'h109b5, 'h107dc, 'h103bc, 'h107ec, 'h109b6, 'h107fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080c, 'h109b7, 'h1081c, 'h1082c, 'h109b8, 'h1083c, 'h1084c, 'h109b9, 'h10bbc, 'h1085c, 'h1086c, 'h109ba, 'h1087c, 'h1088c, 'h109bb, 'h103bc, 'h1089c, 'h108ac, 'h109bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bc, 'h108cc, 'h109bd, 'h108dc, 'h106ec, 'h109be, 'h10bcc, 'h106fc, 'h1070c, 'h109bf, 'h1071c, 'h1072c, 'h109c0, 'h1073c, 'h103bc, 'h1074c, 'h109c1, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076c, 'h109c2, 'h1077c, 'h1078c, 'h109c3, 'h1079c, 'h10bcc, 'h107ac, 'h109c4, 'h107bc, 'h107cc, 'h109c5, 'h107dc, 'h107ec, 'h109c6, 'h103bc, 'h107fc, 'h1080c, 'h109c7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081c, 'h1082c, 'h109c8, 'h1083c, 'h1084c, 'h109c9, 'h10bcc, 'h1085c, 'h1086c, 'h109ca, 'h1087c, 'h1088c, 'h109cb, 'h1089c, 'h103bc, 'h108ac, 'h109cc, 'h108bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cc, 'h109cd, 'h108dc, 'h106ec, 'h109ce, 'h10bdc, 'h106fc, 'h1070c, 'h109cf, 'h1071c, 'h1072c, 'h109d0, 'h1073c, 'h1074c, 'h109d1, 'h103bc, 'h1075c, 'h1076c, 'h109d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077c, 'h1078c, 'h109d3, 'h1079c, 'h10bdc, 'h107ac, 'h109d4, 'h107bc, 'h107cc, 'h109d5, 'h107dc, 'h107ec, 'h109d6, 'h107fc, 'h103bc, 'h1080c, 'h109d7, 'h1081c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082c, 'h109d8, 'h1083c, 'h1084c, 'h109d9, 'h10bdc, 'h1085c, 'h1086c, 'h109da, 'h1087c, 'h1088c, 'h109db, 'h1089c, 'h108ac, 'h109dc, 'h103bc, 'h108bc, 'h108cc, 'h109dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dc, 'h106ec, 'h109de, 'h10bec, 'h106fc, 'h1070c, 'h109df, 'h1071c, 'h1072c, 'h109e0, 'h1073c, 'h1074c, 'h109e1, 'h1075c, 'h103bc, 'h1076c, 'h109e2, 'h1077c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078c, 'h109e3, 'h1079c, 'h10bec, 'h107ac, 'h109e4, 'h107bc, 'h107cc, 'h109e5, 'h107dc, 'h107ec, 'h109e6, 'h107fc, 'h1080c, 'h109e7, 'h103bc, 'h1081c, 'h1082c, 'h109e8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083c, 'h1084c, 'h109e9, 'h10bec, 'h1085c, 'h1086c, 'h109ea, 'h1087c, 'h1088c, 'h109eb, 'h1089c, 'h108ac, 'h109ec, 'h108bc, 'h103bc, 'h108cc, 'h109ed, 'h108dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ec, 'h109ee, 'h10bfc, 'h106fc, 'h1070c, 'h109ef, 'h1071c, 'h1072c, 'h109f0, 'h1073c, 'h1074c, 'h109f1, 'h1075c, 'h1076c, 'h109f2, 'h103bc, 'h1077c, 'h1078c, 'h109f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079c, 'h10bfc, 'h107ac, 'h109f4, 'h107bc, 'h107cc, 'h109f5, 'h107dc, 'h107ec, 'h109f6, 'h107fc, 'h1080c, 'h109f7, 'h1081c, 'h103bc, 'h1082c, 'h109f8, 'h1083c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084c, 'h109f9, 'h10bfc, 'h1085c, 'h1086c, 'h109fa, 'h1087c, 'h1088c, 'h109fb, 'h1089c, 'h108ac, 'h109fc, 'h108bc, 'h108cc, 'h109fd, 'h103bc, 'h108dc, 'h106ec, 'h109fe, 'h10c0c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fc, 'h1070c, 'h109ff, 'h1071c, 'h1072c, 'h10a00, 'h1073c, 'h1074c, 'h10a01, 'h1075c, 'h1076c, 'h10a02, 'h1077c, 'h103bc, 'h1078c, 'h10a03, 'h1079c, 'h10c0c, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ac, 'h10a04, 'h107bc, 'h107cc, 'h10a05, 'h107dc, 'h107ec, 'h10a06, 'h107fc, 'h1080c, 'h10a07, 'h1081c, 'h1082c, 'h10a08, 'h103bc, 'h1083c, 'h1084c, 'h10a09, 'h10c0c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085c, 'h1086c, 'h10a0a, 'h1087c, 'h1088c, 'h10a0b, 'h1089c, 'h108ac, 'h10a0c, 'h108bc, 'h108cc, 'h10a0d, 'h108dc, 'h103bc, 'h106ec, 'h10a0e, 'h10c1c, 'h106fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10a0f, 'h1071c, 'h1072c, 'h10a10, 'h1073c, 'h1074c, 'h10a11, 'h1075c, 'h1076c, 'h10a12, 'h1077c, 'h1078c, 'h10a13, 'h103bc, 'h1079c, 'h10c1c, 'h107ac, 'h10a14, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bc, 'h107cc, 'h10a15, 'h107dc, 'h107ec, 'h10a16, 'h107fc, 'h1080c, 'h10a17, 'h1081c, 'h1082c, 'h10a18, 'h1083c, 'h103bc, 'h1084c, 'h10a19, 'h10c1c, 'h1085c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086c, 'h10a1a, 'h1087c, 'h1088c, 'h10a1b, 'h1089c, 'h108ac, 'h10a1c, 'h108bc, 'h108cc, 'h10a1d, 'h108dc, 'h106ec, 'h10a1e, 'h10c2c, 'h103bc, 'h106fc, 'h1070c, 'h10a1f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071c, 'h1072c, 'h10a20, 'h1073c, 'h1074c, 'h10a21, 'h1075c, 'h1076c, 'h10a22, 'h1077c, 'h1078c, 'h10a23, 'h1079c, 'h10c2c, 'h103bc, 'h107ac, 'h10a24, 'h107bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cc, 'h10a25, 'h107dc, 'h107ec, 'h10a26, 'h107fc, 'h1080c, 'h10a27, 'h1081c, 'h1082c, 'h10a28, 'h1083c, 'h1084c, 'h10a29, 'h10c2c, 'h103bc, 'h1085c, 'h1086c, 'h10a2a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087c, 'h1088c, 'h10a2b, 'h1089c, 'h108ac, 'h10a2c, 'h108bc, 'h108cc, 'h10a2d, 'h108dc, 'h106ec, 'h10a2e, 'h10c3c, 'h106fc, 'h103bc, 'h1070c, 'h10a2f, 'h1071c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072c, 'h10a30, 'h1073c, 'h1074c, 'h10a31, 'h1075c, 'h1076c, 'h10a32, 'h1077c, 'h1078c, 'h10a33, 'h1079c, 'h10c3c, 'h107ac, 'h10a34, 'h103bc, 'h107bc, 'h107cc, 'h10a35, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dc, 'h107ec, 'h10a36, 'h107fc, 'h1080c, 'h10a37, 'h1081c, 'h1082c, 'h10a38, 'h1083c, 'h1084c, 'h10a39, 'h10c3c, 'h1085c, 'h103bc, 'h1086c, 'h10a3a, 'h1087c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088c, 'h10a3b, 'h1089c, 'h108ac, 'h10a3c, 'h108bc, 'h108cc, 'h10a3d, 'h108dc, 'h106ec, 'h10a3e, 'h10c4c, 'h106fc, 'h1070c, 'h10a3f, 'h103bc, 'h1071c, 'h1072c, 'h10a40, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h1074c, 'h10a41, 'h1075c, 'h1076c, 'h10a42, 'h1077c, 'h1078c, 'h10a43, 'h1079c, 'h10c4c, 'h107ac, 'h10a44, 'h107bc, 'h103bc, 'h107cc, 'h10a45, 'h107dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ec, 'h10a46, 'h107fc, 'h1080c, 'h10a47, 'h1081c, 'h1082c, 'h10a48, 'h1083c, 'h1084c, 'h10a49, 'h10c4c, 'h1085c, 'h1086c, 'h10a4a, 'h103bc, 'h1087c, 'h1088c, 'h10a4b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089c, 'h108ac, 'h10a4c, 'h108bc, 'h108cc, 'h10a4d, 'h108dc, 'h106ec, 'h10a4e, 'h10c5c, 'h106fc, 'h1070c, 'h10a4f, 'h1071c, 'h103bc, 'h1072c, 'h10a50, 'h1073c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074c, 'h10a51, 'h1075c, 'h1076c, 'h10a52, 'h1077c, 'h1078c, 'h10a53, 'h1079c, 'h10c5c, 'h107ac, 'h10a54, 'h107bc, 'h107cc, 'h10a55, 'h103bc, 'h107dc, 'h107ec, 'h10a56, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fc, 'h1080c, 'h10a57, 'h1081c, 'h1082c, 'h10a58, 'h1083c, 'h1084c, 'h10a59, 'h10c5c, 'h1085c, 'h1086c, 'h10a5a, 'h1087c, 'h103bc, 'h1088c, 'h10a5b, 'h1089c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ac, 'h10a5c, 'h108bc, 'h108cc, 'h10a5d, 'h108dc, 'h106ec, 'h10a5e, 'h10c6c, 'h106fc, 'h1070c, 'h10a5f, 'h1071c, 'h1072c, 'h10a60, 'h103bc, 'h1073c, 'h1074c, 'h10a61, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075c, 'h1076c, 'h10a62, 'h1077c, 'h1078c, 'h10a63, 'h1079c, 'h10c6c, 'h107ac, 'h10a64, 'h107bc, 'h107cc, 'h10a65, 'h107dc, 'h103bc, 'h107ec, 'h10a66, 'h107fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080c, 'h10a67, 'h1081c, 'h1082c, 'h10a68, 'h1083c, 'h1084c, 'h10a69, 'h10c6c, 'h1085c, 'h1086c, 'h10a6a, 'h1087c, 'h1088c, 'h10a6b, 'h103bc, 'h1089c, 'h108ac, 'h10a6c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bc, 'h108cc, 'h10a6d, 'h108dc, 'h106ec, 'h10a6e, 'h10c7c, 'h106fc, 'h1070c, 'h10a6f, 'h1071c, 'h1072c, 'h10a70, 'h1073c, 'h103bc, 'h1074c, 'h10a71, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076c, 'h10a72, 'h1077c, 'h1078c, 'h10a73, 'h1079c, 'h10c7c, 'h107ac, 'h10a74, 'h107bc, 'h107cc, 'h10a75, 'h107dc, 'h107ec, 'h10a76, 'h103bc, 'h107fc, 'h1080c, 'h10a77, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081c, 'h1082c, 'h10a78, 'h1083c, 'h1084c, 'h10a79, 'h10c7c, 'h1085c, 'h1086c, 'h10a7a, 'h1087c, 'h1088c, 'h10a7b, 'h1089c, 'h103bc, 'h108ac, 'h10a7c, 'h108bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cc, 'h10a7d, 'h108dc, 'h106ec, 'h10a7e, 'h10c8c, 'h106fc, 'h1070c, 'h10a7f, 'h1071c, 'h1072c, 'h10a80, 'h1073c, 'h1074c, 'h10a81, 'h103bc, 'h1075c, 'h1076c, 'h10a82, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077c, 'h1078c, 'h10a83, 'h1079c, 'h10c8c, 'h107ac, 'h10a84, 'h107bc, 'h107cc, 'h10a85, 'h107dc, 'h107ec, 'h10a86, 'h107fc, 'h103bc, 'h1080c, 'h10a87, 'h1081c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082c, 'h10a88, 'h1083c, 'h1084c, 'h10a89, 'h10c8c, 'h1085c, 'h1086c, 'h10a8a, 'h1087c, 'h1088c, 'h10a8b, 'h1089c, 'h108ac, 'h10a8c, 'h103bc, 'h108bc, 'h108cc, 'h10a8d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dc, 'h106ec, 'h10a8e, 'h10c9c, 'h106fc, 'h1070c, 'h10a8f, 'h1071c, 'h1072c, 'h10a90, 'h1073c, 'h1074c, 'h10a91, 'h1075c, 'h103bc, 'h1076c, 'h10a92, 'h1077c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078c, 'h10a93, 'h1079c, 'h10c9c, 'h107ac, 'h10a94, 'h107bc, 'h107cc, 'h10a95, 'h107dc, 'h107ec, 'h10a96, 'h107fc, 'h1080c, 'h10a97, 'h103bc, 'h1081c, 'h1082c, 'h10a98, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083c, 'h1084c, 'h10a99, 'h10c9c, 'h1085c, 'h1086c, 'h10a9a, 'h1087c, 'h1088c, 'h10a9b, 'h1089c, 'h108ac, 'h10a9c, 'h108bc, 'h103bc, 'h108cc, 'h10a9d, 'h108dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ec, 'h10a9e, 'h10cac, 'h106fc, 'h1070c, 'h10a9f, 'h1071c, 'h1072c, 'h10aa0, 'h1073c, 'h1074c, 'h10aa1, 'h1075c, 'h1076c, 'h10aa2, 'h103bc, 'h1077c, 'h1078c, 'h10aa3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079c, 'h10cac, 'h107ac, 'h10aa4, 'h107bc, 'h107cc, 'h10aa5, 'h107dc, 'h107ec, 'h10aa6, 'h107fc, 'h1080c, 'h10aa7, 'h1081c, 'h103bc, 'h1082c, 'h10aa8, 'h1083c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084c, 'h10aa9, 'h10cac, 'h1085c, 'h1086c, 'h10aaa, 'h1087c, 'h1088c, 'h10aab, 'h1089c, 'h108ac, 'h10aac, 'h108bc, 'h108cc, 'h10aad, 'h103bc, 'h108dc, 'h106ec, 'h10aae, 'h10cbc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fc, 'h1070c, 'h10aaf, 'h1071c, 'h1072c, 'h10ab0, 'h1073c, 'h1074c, 'h10ab1, 'h1075c, 'h1076c, 'h10ab2, 'h1077c, 'h103bc, 'h1078c, 'h10ab3, 'h1079c, 'h10cbc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ac, 'h10ab4, 'h107bc, 'h107cc, 'h10ab5, 'h107dc, 'h107ec, 'h10ab6, 'h107fc, 'h1080c, 'h10ab7, 'h1081c, 'h1082c, 'h10ab8, 'h103bc, 'h1083c, 'h1084c, 'h10ab9, 'h10cbc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085c, 'h1086c, 'h10aba, 'h1087c, 'h1088c, 'h10abb, 'h1089c, 'h108ac, 'h10abc, 'h108bc, 'h108cc, 'h10abd, 'h108dc, 'h103bc, 'h106ec, 'h10abe, 'h10ccc, 'h106fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10abf, 'h1071c, 'h1072c, 'h10ac0, 'h1073c, 'h1074c, 'h10ac1, 'h1075c, 'h1076c, 'h10ac2, 'h1077c, 'h1078c, 'h10ac3, 'h103bc, 'h1079c, 'h10ccc, 'h107ac, 'h10ac4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bc, 'h107cc, 'h10ac5, 'h107dc, 'h107ec, 'h10ac6, 'h107fc, 'h1080c, 'h10ac7, 'h1081c, 'h1082c, 'h10ac8, 'h1083c, 'h103bc, 'h1084c, 'h10ac9, 'h10ccc, 'h1085c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086c, 'h10aca, 'h1087c, 'h1088c, 'h10acb, 'h1089c, 'h108ac, 'h10acc, 'h108bc, 'h108cc, 'h10acd, 'h108dc, 'h106ec, 'h10ace, 'h10cdc, 'h103bc, 'h106fc, 'h1070c, 'h10acf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071c, 'h1072c, 'h10ad0, 'h1073c, 'h1074c, 'h10ad1, 'h1075c, 'h1076c, 'h10ad2, 'h1077c, 'h1078c, 'h10ad3, 'h1079c, 'h10cdc, 'h103bc, 'h107ac, 'h10ad4, 'h107bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cc, 'h10ad5, 'h107dc, 'h107ec, 'h10ad6, 'h107fc, 'h1080c, 'h10ad7, 'h1081c, 'h1082c, 'h10ad8, 'h1083c, 'h1084c, 'h10ad9, 'h10cdc, 'h103bc, 'h1085c, 'h1086c, 'h10ada, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087c, 'h1088c, 'h10adb, 'h1089c, 'h108ac, 'h10adc, 'h108bc, 'h108cc, 'h10add, 'h108dc, 'h106ec, 'h108de, 'h10aec, 'h106fc, 'h103bc, 'h1070c, 'h108df, 'h1071c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072c, 'h108e0, 'h1073c, 'h1074c, 'h108e1, 'h1075c, 'h1076c, 'h108e2, 'h1077c, 'h1078c, 'h108e3, 'h1079c, 'h10aec, 'h107ac, 'h108e4, 'h103bc, 'h107bc, 'h107cc, 'h108e5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dc, 'h107ec, 'h108e6, 'h107fc, 'h1080c, 'h108e7, 'h1081c, 'h1082c, 'h108e8, 'h1083c, 'h1084c, 'h108e9, 'h10aec, 'h1085c, 'h103bc, 'h1086c, 'h108ea, 'h1087c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088c, 'h108eb, 'h1089c, 'h108ac, 'h108ec, 'h108bc, 'h108cc, 'h108ed, 'h108dc, 'h106ec, 'h108ee, 'h10afc, 'h106fc, 'h1070c, 'h108ef, 'h103bc, 'h1071c, 'h1072c, 'h108f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h1074c, 'h108f1, 'h1075c, 'h1076c, 'h108f2, 'h1077c, 'h1078c, 'h108f3, 'h1079c, 'h10afc, 'h107ac, 'h108f4, 'h107bc, 'h103bc, 'h107cc, 'h108f5, 'h107dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ec, 'h108f6, 'h107fc, 'h1080c, 'h108f7, 'h1081c, 'h1082c, 'h108f8, 'h1083c, 'h1084c, 'h108f9, 'h10afc, 'h1085c, 'h1086c, 'h108fa, 'h103bc, 'h1087c, 'h1088c, 'h108fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089c, 'h108ac, 'h108fc, 'h108bc, 'h108cc, 'h108fd, 'h108dc, 'h106ec, 'h108fe, 'h10b0c, 'h106fc, 'h1070c, 'h108ff, 'h1071c, 'h103bc, 'h1072c, 'h10900, 'h1073c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074c, 'h10901, 'h1075c, 'h1076c, 'h10902, 'h1077c, 'h1078c, 'h10903, 'h1079c, 'h10b0c, 'h107ac, 'h10904, 'h107bc, 'h107cc, 'h10905, 'h103bc, 'h107dc, 'h107ec, 'h10906, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fc, 'h1080c, 'h10907, 'h1081c, 'h1082c, 'h10908, 'h1083c, 'h1084c, 'h10909, 'h10b0c, 'h1085c, 'h1086c, 'h1090a, 'h1087c, 'h103bc, 'h1088c, 'h1090b, 'h1089c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ac, 'h1090c, 'h108bc, 'h108cc, 'h1090d, 'h108dc, 'h106ec, 'h1090e, 'h10b1c, 'h106fc, 'h1070c, 'h1090f, 'h1071c, 'h1072c, 'h10910, 'h103bc, 'h1073c, 'h1074c, 'h10911, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075c, 'h1076c, 'h10912, 'h1077c, 'h1078c, 'h10913, 'h1079c, 'h10b1c, 'h107ac, 'h10914, 'h107bc, 'h107cc, 'h10915, 'h107dc, 'h103bc, 'h107ec, 'h10916, 'h107fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080c, 'h10917, 'h1081c, 'h1082c, 'h10918, 'h1083c, 'h1084c, 'h10919, 'h10b1c, 'h1085c, 'h1086c, 'h1091a, 'h1087c, 'h1088c, 'h1091b, 'h103bc, 'h1089c, 'h108ac, 'h1091c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bc, 'h108cc, 'h1091d, 'h108dc, 'h106ec, 'h1091e, 'h10b2c, 'h106fc, 'h1070c, 'h1091f, 'h1071c, 'h1072c, 'h10920, 'h1073c, 'h103bc, 'h1074c, 'h10921, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076c, 'h10922, 'h1077c, 'h1078c, 'h10923, 'h1079c, 'h10b2c, 'h107ac, 'h10924, 'h107bc, 'h107cc, 'h10925, 'h107dc, 'h107ec, 'h10926, 'h103bc, 'h107fc, 'h1080c, 'h10927, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081c, 'h1082c, 'h10928, 'h1083c, 'h1084c, 'h10929, 'h10b2c, 'h1085c, 'h1086c, 'h1092a, 'h1087c, 'h1088c, 'h1092b, 'h1089c, 'h103bc, 'h108ac, 'h1092c, 'h108bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cc, 'h1092d, 'h108dc, 'h106ec, 'h1092e, 'h10b3c, 'h106fc, 'h1070c, 'h1092f, 'h1071c, 'h1072c, 'h10930, 'h1073c, 'h1074c, 'h10931, 'h103bc, 'h1075c, 'h1076c, 'h10932, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077c, 'h1078c, 'h10933, 'h1079c, 'h10b3c, 'h107ac, 'h10934, 'h107bc, 'h107cc, 'h10935, 'h107dc, 'h107ec, 'h10936, 'h107fc, 'h103bc, 'h1080c, 'h10937, 'h1081c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082c, 'h10938, 'h1083c, 'h1084c, 'h10939, 'h10b3c, 'h1085c, 'h1086c, 'h1093a, 'h1087c, 'h1088c, 'h1093b, 'h1089c, 'h108ac, 'h1093c, 'h103bc, 'h108bc, 'h108cc, 'h1093d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dc, 'h106ec, 'h1093e, 'h10b4c, 'h106fc, 'h1070c, 'h1093f, 'h1071c, 'h1072c, 'h10940, 'h1073c, 'h1074c, 'h10941, 'h1075c, 'h103bc, 'h1076c, 'h10942, 'h1077c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078c, 'h10943, 'h1079c, 'h10b4c, 'h107ac, 'h10944, 'h107bc, 'h107cc, 'h10945, 'h107dc, 'h107ec, 'h10946, 'h107fc, 'h1080c, 'h10947, 'h103bc, 'h1081c, 'h1082c, 'h10948, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083c, 'h1084c, 'h10949, 'h10b4c, 'h1085c, 'h1086c, 'h1094a, 'h1087c, 'h1088c, 'h1094b, 'h1089c, 'h108ac, 'h1094c, 'h108bc, 'h103bc, 'h108cc, 'h1094d, 'h108dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ec, 'h1094e, 'h10b5c, 'h106fc, 'h1070c, 'h1094f, 'h1071c, 'h1072c, 'h10950, 'h1073c, 'h1074c, 'h10951, 'h1075c, 'h1076c, 'h10952, 'h103bc, 'h1077c, 'h1078c, 'h10953, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079c, 'h10b5c, 'h107ac, 'h10954, 'h107bc, 'h107cc, 'h10955, 'h107dc, 'h107ec, 'h10956, 'h107fc, 'h1080c, 'h10957, 'h1081c, 'h103bc, 'h1082c, 'h10958, 'h1083c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084c, 'h10959, 'h10b5c, 'h1085c, 'h1086c, 'h1095a, 'h1087c, 'h1088c, 'h1095b, 'h1089c, 'h108ac, 'h1095c, 'h108bc, 'h108cc, 'h1095d, 'h103bc, 'h108dc, 'h106ec, 'h1095e, 'h10b6c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fc, 'h1070c, 'h1095f, 'h1071c, 'h1072c, 'h10960, 'h1073c, 'h1074c, 'h10961, 'h1075c, 'h1076c, 'h10962, 'h1077c, 'h103bc, 'h1078c, 'h10963, 'h1079c, 'h10b6c, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ac, 'h10964, 'h107bc, 'h107cc, 'h10965, 'h107dc, 'h107ec, 'h10966, 'h107fc, 'h1080c, 'h10967, 'h1081c, 'h1082c, 'h10968, 'h103bc, 'h1083c, 'h1084c, 'h10969, 'h10b6c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085c, 'h1086c, 'h1096a, 'h1087c, 'h1088c, 'h1096b, 'h1089c, 'h108ac, 'h1096c, 'h108bc, 'h108cc, 'h1096d, 'h108dc, 'h103bc, 'h106ec, 'h1096e, 'h10b7c, 'h106fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h1096f, 'h1071c, 'h1072c, 'h10970, 'h1073c, 'h1074c, 'h10971, 'h1075c, 'h1076c, 'h10972, 'h1077c, 'h1078c, 'h10973, 'h103bc, 'h1079c, 'h10b7c, 'h107ac, 'h10974, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bc, 'h107cc, 'h10975, 'h107dc, 'h107ec, 'h10976, 'h107fc, 'h1080c, 'h10977, 'h1081c, 'h1082c, 'h10978, 'h1083c, 'h103bc, 'h1084c, 'h10979, 'h10b7c, 'h1085c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086c, 'h1097a, 'h1087c, 'h1088c, 'h1097b, 'h1089c, 'h108ac, 'h1097c, 'h108bc, 'h108cc, 'h1097d, 'h108dc, 'h106ec, 'h1097e, 'h10b8c, 'h103bc, 'h106fc, 'h1070c, 'h1097f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071c, 'h1072c, 'h10980, 'h1073c, 'h1074c, 'h10981, 'h1075c, 'h1076c, 'h10982, 'h1077c, 'h1078c, 'h10983, 'h1079c, 'h10b8c, 'h103bc, 'h107ac, 'h10984, 'h107bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cc, 'h10985, 'h107dc, 'h107ec, 'h10986, 'h107fc, 'h1080c, 'h10987, 'h1081c, 'h1082c, 'h10988, 'h1083c, 'h1084c, 'h10989, 'h10b8c, 'h103bc, 'h1085c, 'h1086c, 'h1098a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087c, 'h1088c, 'h1098b, 'h1089c, 'h108ac, 'h1098c, 'h108bc, 'h108cc, 'h1098d, 'h108dc, 'h106ec, 'h1098e, 'h10b9c, 'h106fc, 'h103bc, 'h1070c, 'h1098f, 'h1071c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072c, 'h10990, 'h1073c, 'h1074c, 'h10991, 'h1075c, 'h1076c, 'h10992, 'h1077c, 'h1078c, 'h10993, 'h1079c, 'h10b9c, 'h107ac, 'h10994, 'h103bc, 'h107bc, 'h107cc, 'h10995, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dc, 'h107ec, 'h10996, 'h107fc, 'h1080c, 'h10997, 'h1081c, 'h1082c, 'h10998, 'h1083c, 'h1084c, 'h10999, 'h10b9c, 'h1085c, 'h103bc, 'h1086c, 'h1099a, 'h1087c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088c, 'h1099b, 'h1089c, 'h108ac, 'h1099c, 'h108bc, 'h108cc, 'h1099d, 'h108dc, 'h106ec, 'h1099e, 'h10bac, 'h106fc, 'h1070c, 'h1099f, 'h103bc, 'h1071c, 'h1072c, 'h109a0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h1074c, 'h109a1, 'h1075c, 'h1076c, 'h109a2, 'h1077c, 'h1078c, 'h109a3, 'h1079c, 'h10bac, 'h107ac, 'h109a4, 'h107bc, 'h103bc, 'h107cc, 'h109a5, 'h107dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ec, 'h109a6, 'h107fc, 'h1080c, 'h109a7, 'h1081c, 'h1082c, 'h109a8, 'h1083c, 'h1084c, 'h109a9, 'h10bac, 'h1085c, 'h1086c, 'h109aa, 'h103bc, 'h1087c, 'h1088c, 'h109ab, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089c, 'h108ac, 'h109ac, 'h108bc, 'h108cc, 'h109ad, 'h108dc, 'h106ec, 'h109ae, 'h10bbc, 'h106fc, 'h1070c, 'h109af, 'h1071c, 'h103bc, 'h1072c, 'h109b0, 'h1073c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074c, 'h109b1, 'h1075c, 'h1076c, 'h109b2, 'h1077c, 'h1078c, 'h109b3, 'h1079c, 'h10bbc, 'h107ac, 'h109b4, 'h107bc, 'h107cc, 'h109b5, 'h103bc, 'h107dc, 'h107ec, 'h109b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fc, 'h1080c, 'h109b7, 'h1081c, 'h1082c, 'h109b8, 'h1083c, 'h1084c, 'h109b9, 'h10bbc, 'h1085c, 'h1086c, 'h109ba, 'h1087c, 'h103bc, 'h1088c, 'h109bb, 'h1089c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ac, 'h109bc, 'h108bc, 'h108cc, 'h109bd, 'h108dc, 'h106ec, 'h109be, 'h10bcc, 'h106fc, 'h1070c, 'h109bf, 'h1071c, 'h1072c, 'h109c0, 'h103bc, 'h1073c, 'h1074c, 'h109c1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075c, 'h1076c, 'h109c2, 'h1077c, 'h1078c, 'h109c3, 'h1079c, 'h10bcc, 'h107ac, 'h109c4, 'h107bc, 'h107cc, 'h109c5, 'h107dc, 'h103bc, 'h107ec, 'h109c6, 'h107fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080c, 'h109c7, 'h1081c, 'h1082c, 'h109c8, 'h1083c, 'h1084c, 'h109c9, 'h10bcc, 'h1085c, 'h1086c, 'h109ca, 'h1087c, 'h1088c, 'h109cb, 'h103bc, 'h1089c, 'h108ac, 'h109cc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bc, 'h108cc, 'h109cd, 'h108dc, 'h106ec, 'h109ce, 'h10bdc, 'h106fc, 'h1070c, 'h109cf, 'h1071c, 'h1072c, 'h109d0, 'h1073c, 'h103bc, 'h1074c, 'h109d1, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076c, 'h109d2, 'h1077c, 'h1078c, 'h109d3, 'h1079c, 'h10bdc, 'h107ac, 'h109d4, 'h107bc, 'h107cc, 'h109d5, 'h107dc, 'h107ec, 'h109d6, 'h103bc, 'h107fc, 'h1080c, 'h109d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081c, 'h1082c, 'h109d8, 'h1083c, 'h1084c, 'h109d9, 'h10bdc, 'h1085c, 'h1086c, 'h109da, 'h1087c, 'h1088c, 'h109db, 'h1089c, 'h103bc, 'h108ac, 'h109dc, 'h108bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cc, 'h109dd, 'h108dc, 'h106ec, 'h109de, 'h10bec, 'h106fc, 'h1070c, 'h109df, 'h1071c, 'h1072c, 'h109e0, 'h1073c, 'h1074c, 'h109e1, 'h103bc, 'h1075c, 'h1076c, 'h109e2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077c, 'h1078c, 'h109e3, 'h1079c, 'h10bec, 'h107ac, 'h109e4, 'h107bc, 'h107cc, 'h109e5, 'h107dc, 'h107ec, 'h109e6, 'h107fc, 'h103bc, 'h1080c, 'h109e7, 'h1081c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082c, 'h109e8, 'h1083c, 'h1084c, 'h109e9, 'h10bec, 'h1085c, 'h1086c, 'h109ea, 'h1087c, 'h1088c, 'h109eb, 'h1089c, 'h108ac, 'h109ec, 'h103bc, 'h108bc, 'h108cc, 'h109ed, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dc, 'h106ec, 'h109ee, 'h10bfc, 'h106fc, 'h1070c, 'h109ef, 'h1071c, 'h1072c, 'h109f0, 'h1073c, 'h1074c, 'h109f1, 'h1075c, 'h103bc, 'h1076c, 'h109f2, 'h1077c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078c, 'h109f3, 'h1079c, 'h10bfc, 'h107ac, 'h109f4, 'h107bc, 'h107cc, 'h109f5, 'h107dc, 'h107ec, 'h109f6, 'h107fc, 'h1080c, 'h109f7, 'h103bc, 'h1081c, 'h1082c, 'h109f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083c, 'h1084c, 'h109f9, 'h10bfc, 'h1085c, 'h1086c, 'h109fa, 'h1087c, 'h1088c, 'h109fb, 'h1089c, 'h108ac, 'h109fc, 'h108bc, 'h103bc, 'h108cc, 'h109fd, 'h108dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ec, 'h109fe, 'h10c0c, 'h106fc, 'h1070c, 'h109ff, 'h1071c, 'h1072c, 'h10a00, 'h1073c, 'h1074c, 'h10a01, 'h1075c, 'h1076c, 'h10a02, 'h103bc, 'h1077c, 'h1078c, 'h10a03, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079c, 'h10c0c, 'h107ac, 'h10a04, 'h107bc, 'h107cc, 'h10a05, 'h107dc, 'h107ec, 'h10a06, 'h107fc, 'h1080c, 'h10a07, 'h1081c, 'h103bc, 'h1082c, 'h10a08, 'h1083c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084c, 'h10a09, 'h10c0c, 'h1085c, 'h1086c, 'h10a0a, 'h1087c, 'h1088c, 'h10a0b, 'h1089c, 'h108ac, 'h10a0c, 'h108bc, 'h108cc, 'h10a0d, 'h103bc, 'h108dc, 'h106ec, 'h10a0e, 'h10c1c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fc, 'h1070c, 'h10a0f, 'h1071c, 'h1072c, 'h10a10, 'h1073c, 'h1074c, 'h10a11, 'h1075c, 'h1076c, 'h10a12, 'h1077c, 'h103bc, 'h1078c, 'h10a13, 'h1079c, 'h10c1c, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ac, 'h10a14, 'h107bc, 'h107cc, 'h10a15, 'h107dc, 'h107ec, 'h10a16, 'h107fc, 'h1080c, 'h10a17, 'h1081c, 'h1082c, 'h10a18, 'h103bc, 'h1083c, 'h1084c, 'h10a19, 'h10c1c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085c, 'h1086c, 'h10a1a, 'h1087c, 'h1088c, 'h10a1b, 'h1089c, 'h108ac, 'h10a1c, 'h108bc, 'h108cc, 'h10a1d, 'h108dc, 'h103bc, 'h106ec, 'h10a1e, 'h10c2c, 'h106fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10a1f, 'h1071c, 'h1072c, 'h10a20, 'h1073c, 'h1074c, 'h10a21, 'h1075c, 'h1076c, 'h10a22, 'h1077c, 'h1078c, 'h10a23, 'h103bc, 'h1079c, 'h10c2c, 'h107ac, 'h10a24, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bc, 'h107cc, 'h10a25, 'h107dc, 'h107ec, 'h10a26, 'h107fc, 'h1080c, 'h10a27, 'h1081c, 'h1082c, 'h10a28, 'h1083c, 'h103bc, 'h1084c, 'h10a29, 'h10c2c, 'h1085c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086c, 'h10a2a, 'h1087c, 'h1088c, 'h10a2b, 'h1089c, 'h108ac, 'h10a2c, 'h108bc, 'h108cc, 'h10a2d, 'h108dc, 'h106ec, 'h10a2e, 'h10c3c, 'h103bc, 'h106fc, 'h1070c, 'h10a2f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071c, 'h1072c, 'h10a30, 'h1073c, 'h1074c, 'h10a31, 'h1075c, 'h1076c, 'h10a32, 'h1077c, 'h1078c, 'h10a33, 'h1079c, 'h10c3c, 'h103bc, 'h107ac, 'h10a34, 'h107bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cc, 'h10a35, 'h107dc, 'h107ec, 'h10a36, 'h107fc, 'h1080c, 'h10a37, 'h1081c, 'h1082c, 'h10a38, 'h1083c, 'h1084c, 'h10a39, 'h10c3c, 'h103bc, 'h1085c, 'h1086c, 'h10a3a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087c, 'h1088c, 'h10a3b, 'h1089c, 'h108ac, 'h10a3c, 'h108bc, 'h108cc, 'h10a3d, 'h108dc, 'h106ec, 'h10a3e, 'h10c4c, 'h106fc, 'h103bc, 'h1070c, 'h10a3f, 'h1071c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072c, 'h10a40, 'h1073c, 'h1074c, 'h10a41, 'h1075c, 'h1076c, 'h10a42, 'h1077c, 'h1078c, 'h10a43, 'h1079c, 'h10c4c, 'h107ac, 'h10a44, 'h103bc, 'h107bc, 'h107cc, 'h10a45, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dc, 'h107ec, 'h10a46, 'h107fc, 'h1080c, 'h10a47, 'h1081c, 'h1082c, 'h10a48, 'h1083c, 'h1084c, 'h10a49, 'h10c4c, 'h1085c, 'h103bc, 'h1086c, 'h10a4a, 'h1087c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088c, 'h10a4b, 'h1089c, 'h108ac, 'h10a4c, 'h108bc, 'h108cc, 'h10a4d, 'h108dc, 'h106ec, 'h10a4e, 'h10c5c, 'h106fc, 'h1070c, 'h10a4f, 'h103bc, 'h1071c, 'h1072c, 'h10a50, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h1074c, 'h10a51, 'h1075c, 'h1076c, 'h10a52, 'h1077c, 'h1078c, 'h10a53, 'h1079c, 'h10c5c, 'h107ac, 'h10a54, 'h107bc, 'h103bc, 'h107cc, 'h10a55, 'h107dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ec, 'h10a56, 'h107fc, 'h1080c, 'h10a57, 'h1081c, 'h1082c, 'h10a58, 'h1083c, 'h1084c, 'h10a59, 'h10c5c, 'h1085c, 'h1086c, 'h10a5a, 'h103bc, 'h1087c, 'h1088c, 'h10a5b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089c, 'h108ac, 'h10a5c, 'h108bc, 'h108cc, 'h10a5d, 'h108dc, 'h106ec, 'h10a5e, 'h10c6c, 'h106fc, 'h1070c, 'h10a5f, 'h1071c, 'h103bc, 'h1072c, 'h10a60, 'h1073c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074c, 'h10a61, 'h1075c, 'h1076c, 'h10a62, 'h1077c, 'h1078c, 'h10a63, 'h1079c, 'h10c6c, 'h107ac, 'h10a64, 'h107bc, 'h107cc, 'h10a65, 'h103bc, 'h107dc, 'h107ec, 'h10a66, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fc, 'h1080c, 'h10a67, 'h1081c, 'h1082c, 'h10a68, 'h1083c, 'h1084c, 'h10a69, 'h10c6c, 'h1085c, 'h1086c, 'h10a6a, 'h1087c, 'h103bc, 'h1088c, 'h10a6b, 'h1089c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ac, 'h10a6c, 'h108bc, 'h108cc, 'h10a6d, 'h108dc, 'h106ec, 'h10a6e, 'h10c7c, 'h106fc, 'h1070c, 'h10a6f, 'h1071c, 'h1072c, 'h10a70, 'h103bc, 'h1073c, 'h1074c, 'h10a71, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075c, 'h1076c, 'h10a72, 'h1077c, 'h1078c, 'h10a73, 'h1079c, 'h10c7c, 'h107ac, 'h10a74, 'h107bc, 'h107cc, 'h10a75, 'h107dc, 'h103bc, 'h107ec, 'h10a76, 'h107fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080c, 'h10a77, 'h1081c, 'h1082c, 'h10a78, 'h1083c, 'h1084c, 'h10a79, 'h10c7c, 'h1085c, 'h1086c, 'h10a7a, 'h1087c, 'h1088c, 'h10a7b, 'h103bc, 'h1089c, 'h108ac, 'h10a7c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bc, 'h108cc, 'h10a7d, 'h108dc, 'h106ec, 'h10a7e, 'h10c8c, 'h106fc, 'h1070c, 'h10a7f, 'h1071c, 'h1072c, 'h10a80, 'h1073c, 'h103bc, 'h1074c, 'h10a81, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076c, 'h10a82, 'h1077c, 'h1078c, 'h10a83, 'h1079c, 'h10c8c, 'h107ac, 'h10a84, 'h107bc, 'h107cc, 'h10a85, 'h107dc, 'h107ec, 'h10a86, 'h103bc, 'h107fc, 'h1080c, 'h10a87, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081c, 'h1082c, 'h10a88, 'h1083c, 'h1084c, 'h10a89, 'h10c8c, 'h1085c, 'h1086c, 'h10a8a, 'h1087c, 'h1088c, 'h10a8b, 'h1089c, 'h103bc, 'h108ac, 'h10a8c, 'h108bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cc, 'h10a8d, 'h108dc, 'h106ec, 'h10a8e, 'h10c9c, 'h106fc, 'h1070c, 'h10a8f, 'h1071c, 'h1072c, 'h10a90, 'h1073c, 'h1074c, 'h10a91, 'h103bc, 'h1075c, 'h1076c, 'h10a92, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077c, 'h1078c, 'h10a93, 'h1079c, 'h10c9c, 'h107ac, 'h10a94, 'h107bc, 'h107cc, 'h10a95, 'h107dc, 'h107ec, 'h10a96, 'h107fc, 'h103bc, 'h1080c, 'h10a97, 'h1081c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082c, 'h10a98, 'h1083c, 'h1084c, 'h10a99, 'h10c9c, 'h1085c, 'h1086c, 'h10a9a, 'h1087c, 'h1088c, 'h10a9b, 'h1089c, 'h108ac, 'h10a9c, 'h103bc, 'h108bc, 'h108cc, 'h10a9d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dc, 'h106ec, 'h10a9e, 'h10cac, 'h106fc, 'h1070c, 'h10a9f, 'h1071c, 'h1072c, 'h10aa0, 'h1073c, 'h1074c, 'h10aa1, 'h1075c, 'h103bc, 'h1076c, 'h10aa2, 'h1077c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078c, 'h10aa3, 'h1079c, 'h10cac, 'h107ac, 'h10aa4, 'h107bc, 'h107cc, 'h10aa5, 'h107dc, 'h107ec, 'h10aa6, 'h107fc, 'h1080c, 'h10aa7, 'h103bc, 'h1081c, 'h1082c, 'h10aa8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083c, 'h1084c, 'h10aa9, 'h10cac, 'h1085c, 'h1086c, 'h10aaa, 'h1087c, 'h1088c, 'h10aab, 'h1089c, 'h108ac, 'h10aac, 'h108bc, 'h103bc, 'h108cc, 'h10aad, 'h108dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ec, 'h10aae, 'h10cbc, 'h106fc, 'h1070c, 'h10aaf, 'h1071c, 'h1072c, 'h10ab0, 'h1073c, 'h1074c, 'h10ab1, 'h1075c, 'h1076c, 'h10ab2, 'h103bc, 'h1077c, 'h1078c, 'h10ab3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079c, 'h10cbc, 'h107ac, 'h10ab4, 'h107bc, 'h107cc, 'h10ab5, 'h107dc, 'h107ec, 'h10ab6, 'h107fc, 'h1080c, 'h10ab7, 'h1081c, 'h103bc, 'h1082c, 'h10ab8, 'h1083c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084c, 'h10ab9, 'h10cbc, 'h1085c, 'h1086c, 'h10aba, 'h1087c, 'h1088c, 'h10abb, 'h1089c, 'h108ac, 'h10abc, 'h108bc, 'h108cc, 'h10abd, 'h103bc, 'h108dc, 'h106ec, 'h10abe, 'h10ccc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fc, 'h1070c, 'h10abf, 'h1071c, 'h1072c, 'h10ac0, 'h1073c, 'h1074c, 'h10ac1, 'h1075c, 'h1076c, 'h10ac2, 'h1077c, 'h103bc, 'h1078c, 'h10ac3, 'h1079c, 'h10ccc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ac, 'h10ac4, 'h107bc, 'h107cc, 'h10ac5, 'h107dc, 'h107ec, 'h10ac6, 'h107fc, 'h1080c, 'h10ac7, 'h1081c, 'h1082c, 'h10ac8, 'h103bc, 'h1083c, 'h1084c, 'h10ac9, 'h10ccc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085c, 'h1086c, 'h10aca, 'h1087c, 'h1088c, 'h10acb, 'h1089c, 'h108ac, 'h10acc, 'h108bc, 'h108cc, 'h10acd, 'h108dc, 'h103bc, 'h106ec, 'h10ace, 'h10cdc, 'h106fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10acf, 'h1071c, 'h1072c, 'h10ad0, 'h1073c, 'h1074c, 'h10ad1, 'h1075c, 'h1076c, 'h10ad2, 'h1077c, 'h1078c, 'h10ad3, 'h103bc, 'h1079c, 'h10cdc, 'h107ac, 'h10ad4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bc, 'h107cc, 'h10ad5, 'h107dc, 'h107ec, 'h10ad6, 'h107fc, 'h1080c, 'h10ad7, 'h1081c, 'h1082c, 'h10ad8, 'h1083c, 'h103bc, 'h1084c, 'h10ad9, 'h10cdc, 'h1085c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086c, 'h10ada, 'h1087c, 'h1088c, 'h10adb, 'h1089c, 'h108ac, 'h10adc, 'h108bc, 'h108cc, 'h10add, 'h108dc, 'h106ed, 'h108de, 'h10aed, 'h103bc, 'h106fd, 'h1070d, 'h108df, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071d, 'h1072d, 'h108e0, 'h1073d, 'h1074d, 'h108e1, 'h1075d, 'h1076d, 'h108e2, 'h1077d, 'h1078d, 'h108e3, 'h1079d, 'h10aed, 'h103bc, 'h107ad, 'h108e4, 'h107bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cd, 'h108e5, 'h107dd, 'h107ed, 'h108e6, 'h107fd, 'h1080d, 'h108e7, 'h1081d, 'h1082d, 'h108e8, 'h1083d, 'h1084d, 'h108e9, 'h10aed, 'h103bc, 'h1085d, 'h1086d, 'h108ea, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087d, 'h1088d, 'h108eb, 'h1089d, 'h108ad, 'h108ec, 'h108bd, 'h108cd, 'h108ed, 'h108dd, 'h106ed, 'h108ee, 'h10afd, 'h106fd, 'h103bc, 'h1070d, 'h108ef, 'h1071d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072d, 'h108f0, 'h1073d, 'h1074d, 'h108f1, 'h1075d, 'h1076d, 'h108f2, 'h1077d, 'h1078d, 'h108f3, 'h1079d, 'h10afd, 'h107ad, 'h108f4, 'h103bc, 'h107bd, 'h107cd, 'h108f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dd, 'h107ed, 'h108f6, 'h107fd, 'h1080d, 'h108f7, 'h1081d, 'h1082d, 'h108f8, 'h1083d, 'h1084d, 'h108f9, 'h10afd, 'h1085d, 'h103bc, 'h1086d, 'h108fa, 'h1087d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088d, 'h108fb, 'h1089d, 'h108ad, 'h108fc, 'h108bd, 'h108cd, 'h108fd, 'h108dd, 'h106ed, 'h108fe, 'h10b0d, 'h106fd, 'h1070d, 'h108ff, 'h103bc, 'h1071d, 'h1072d, 'h10900, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h1074d, 'h10901, 'h1075d, 'h1076d, 'h10902, 'h1077d, 'h1078d, 'h10903, 'h1079d, 'h10b0d, 'h107ad, 'h10904, 'h107bd, 'h103bc, 'h107cd, 'h10905, 'h107dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ed, 'h10906, 'h107fd, 'h1080d, 'h10907, 'h1081d, 'h1082d, 'h10908, 'h1083d, 'h1084d, 'h10909, 'h10b0d, 'h1085d, 'h1086d, 'h1090a, 'h103bc, 'h1087d, 'h1088d, 'h1090b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089d, 'h108ad, 'h1090c, 'h108bd, 'h108cd, 'h1090d, 'h108dd, 'h106ed, 'h1090e, 'h10b1d, 'h106fd, 'h1070d, 'h1090f, 'h1071d, 'h103bc, 'h1072d, 'h10910, 'h1073d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074d, 'h10911, 'h1075d, 'h1076d, 'h10912, 'h1077d, 'h1078d, 'h10913, 'h1079d, 'h10b1d, 'h107ad, 'h10914, 'h107bd, 'h107cd, 'h10915, 'h103bc, 'h107dd, 'h107ed, 'h10916, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fd, 'h1080d, 'h10917, 'h1081d, 'h1082d, 'h10918, 'h1083d, 'h1084d, 'h10919, 'h10b1d, 'h1085d, 'h1086d, 'h1091a, 'h1087d, 'h103bc, 'h1088d, 'h1091b, 'h1089d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ad, 'h1091c, 'h108bd, 'h108cd, 'h1091d, 'h108dd, 'h106ed, 'h1091e, 'h10b2d, 'h106fd, 'h1070d, 'h1091f, 'h1071d, 'h1072d, 'h10920, 'h103bc, 'h1073d, 'h1074d, 'h10921, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075d, 'h1076d, 'h10922, 'h1077d, 'h1078d, 'h10923, 'h1079d, 'h10b2d, 'h107ad, 'h10924, 'h107bd, 'h107cd, 'h10925, 'h107dd, 'h103bc, 'h107ed, 'h10926, 'h107fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080d, 'h10927, 'h1081d, 'h1082d, 'h10928, 'h1083d, 'h1084d, 'h10929, 'h10b2d, 'h1085d, 'h1086d, 'h1092a, 'h1087d, 'h1088d, 'h1092b, 'h103bc, 'h1089d, 'h108ad, 'h1092c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bd, 'h108cd, 'h1092d, 'h108dd, 'h106ed, 'h1092e, 'h10b3d, 'h106fd, 'h1070d, 'h1092f, 'h1071d, 'h1072d, 'h10930, 'h1073d, 'h103bc, 'h1074d, 'h10931, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076d, 'h10932, 'h1077d, 'h1078d, 'h10933, 'h1079d, 'h10b3d, 'h107ad, 'h10934, 'h107bd, 'h107cd, 'h10935, 'h107dd, 'h107ed, 'h10936, 'h103bc, 'h107fd, 'h1080d, 'h10937, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081d, 'h1082d, 'h10938, 'h1083d, 'h1084d, 'h10939, 'h10b3d, 'h1085d, 'h1086d, 'h1093a, 'h1087d, 'h1088d, 'h1093b, 'h1089d, 'h103bc, 'h108ad, 'h1093c, 'h108bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cd, 'h1093d, 'h108dd, 'h106ed, 'h1093e, 'h10b4d, 'h106fd, 'h1070d, 'h1093f, 'h1071d, 'h1072d, 'h10940, 'h1073d, 'h1074d, 'h10941, 'h103bc, 'h1075d, 'h1076d, 'h10942, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077d, 'h1078d, 'h10943, 'h1079d, 'h10b4d, 'h107ad, 'h10944, 'h107bd, 'h107cd, 'h10945, 'h107dd, 'h107ed, 'h10946, 'h107fd, 'h103bc, 'h1080d, 'h10947, 'h1081d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082d, 'h10948, 'h1083d, 'h1084d, 'h10949, 'h10b4d, 'h1085d, 'h1086d, 'h1094a, 'h1087d, 'h1088d, 'h1094b, 'h1089d, 'h108ad, 'h1094c, 'h103bc, 'h108bd, 'h108cd, 'h1094d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dd, 'h106ed, 'h1094e, 'h10b5d, 'h106fd, 'h1070d, 'h1094f, 'h1071d, 'h1072d, 'h10950, 'h1073d, 'h1074d, 'h10951, 'h1075d, 'h103bc, 'h1076d, 'h10952, 'h1077d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078d, 'h10953, 'h1079d, 'h10b5d, 'h107ad, 'h10954, 'h107bd, 'h107cd, 'h10955, 'h107dd, 'h107ed, 'h10956, 'h107fd, 'h1080d, 'h10957, 'h103bc, 'h1081d, 'h1082d, 'h10958, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083d, 'h1084d, 'h10959, 'h10b5d, 'h1085d, 'h1086d, 'h1095a, 'h1087d, 'h1088d, 'h1095b, 'h1089d, 'h108ad, 'h1095c, 'h108bd, 'h103bc, 'h108cd, 'h1095d, 'h108dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ed, 'h1095e, 'h10b6d, 'h106fd, 'h1070d, 'h1095f, 'h1071d, 'h1072d, 'h10960, 'h1073d, 'h1074d, 'h10961, 'h1075d, 'h1076d, 'h10962, 'h103bc, 'h1077d, 'h1078d, 'h10963, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079d, 'h10b6d, 'h107ad, 'h10964, 'h107bd, 'h107cd, 'h10965, 'h107dd, 'h107ed, 'h10966, 'h107fd, 'h1080d, 'h10967, 'h1081d, 'h103bc, 'h1082d, 'h10968, 'h1083d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084d, 'h10969, 'h10b6d, 'h1085d, 'h1086d, 'h1096a, 'h1087d, 'h1088d, 'h1096b, 'h1089d, 'h108ad, 'h1096c, 'h108bd, 'h108cd, 'h1096d, 'h103bc, 'h108dd, 'h106ed, 'h1096e, 'h10b7d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fd, 'h1070d, 'h1096f, 'h1071d, 'h1072d, 'h10970, 'h1073d, 'h1074d, 'h10971, 'h1075d, 'h1076d, 'h10972, 'h1077d, 'h103bc, 'h1078d, 'h10973, 'h1079d, 'h10b7d, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ad, 'h10974, 'h107bd, 'h107cd, 'h10975, 'h107dd, 'h107ed, 'h10976, 'h107fd, 'h1080d, 'h10977, 'h1081d, 'h1082d, 'h10978, 'h103bc, 'h1083d, 'h1084d, 'h10979, 'h10b7d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085d, 'h1086d, 'h1097a, 'h1087d, 'h1088d, 'h1097b, 'h1089d, 'h108ad, 'h1097c, 'h108bd, 'h108cd, 'h1097d, 'h108dd, 'h103bc, 'h106ed, 'h1097e, 'h10b8d, 'h106fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h1097f, 'h1071d, 'h1072d, 'h10980, 'h1073d, 'h1074d, 'h10981, 'h1075d, 'h1076d, 'h10982, 'h1077d, 'h1078d, 'h10983, 'h103bc, 'h1079d, 'h10b8d, 'h107ad, 'h10984, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bd, 'h107cd, 'h10985, 'h107dd, 'h107ed, 'h10986, 'h107fd, 'h1080d, 'h10987, 'h1081d, 'h1082d, 'h10988, 'h1083d, 'h103bc, 'h1084d, 'h10989, 'h10b8d, 'h1085d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086d, 'h1098a, 'h1087d, 'h1088d, 'h1098b, 'h1089d, 'h108ad, 'h1098c, 'h108bd, 'h108cd, 'h1098d, 'h108dd, 'h106ed, 'h1098e, 'h10b9d, 'h103bc, 'h106fd, 'h1070d, 'h1098f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071d, 'h1072d, 'h10990, 'h1073d, 'h1074d, 'h10991, 'h1075d, 'h1076d, 'h10992, 'h1077d, 'h1078d, 'h10993, 'h1079d, 'h10b9d, 'h103bc, 'h107ad, 'h10994, 'h107bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cd, 'h10995, 'h107dd, 'h107ed, 'h10996, 'h107fd, 'h1080d, 'h10997, 'h1081d, 'h1082d, 'h10998, 'h1083d, 'h1084d, 'h10999, 'h10b9d, 'h103bc, 'h1085d, 'h1086d, 'h1099a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087d, 'h1088d, 'h1099b, 'h1089d, 'h108ad, 'h1099c, 'h108bd, 'h108cd, 'h1099d, 'h108dd, 'h106ed, 'h1099e, 'h10bad, 'h106fd, 'h103bc, 'h1070d, 'h1099f, 'h1071d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072d, 'h109a0, 'h1073d, 'h1074d, 'h109a1, 'h1075d, 'h1076d, 'h109a2, 'h1077d, 'h1078d, 'h109a3, 'h1079d, 'h10bad, 'h107ad, 'h109a4, 'h103bc, 'h107bd, 'h107cd, 'h109a5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dd, 'h107ed, 'h109a6, 'h107fd, 'h1080d, 'h109a7, 'h1081d, 'h1082d, 'h109a8, 'h1083d, 'h1084d, 'h109a9, 'h10bad, 'h1085d, 'h103bc, 'h1086d, 'h109aa, 'h1087d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088d, 'h109ab, 'h1089d, 'h108ad, 'h109ac, 'h108bd, 'h108cd, 'h109ad, 'h108dd, 'h106ed, 'h109ae, 'h10bbd, 'h106fd, 'h1070d, 'h109af, 'h103bc, 'h1071d, 'h1072d, 'h109b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h1074d, 'h109b1, 'h1075d, 'h1076d, 'h109b2, 'h1077d, 'h1078d, 'h109b3, 'h1079d, 'h10bbd, 'h107ad, 'h109b4, 'h107bd, 'h103bc, 'h107cd, 'h109b5, 'h107dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ed, 'h109b6, 'h107fd, 'h1080d, 'h109b7, 'h1081d, 'h1082d, 'h109b8, 'h1083d, 'h1084d, 'h109b9, 'h10bbd, 'h1085d, 'h1086d, 'h109ba, 'h103bc, 'h1087d, 'h1088d, 'h109bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089d, 'h108ad, 'h109bc, 'h108bd, 'h108cd, 'h109bd, 'h108dd, 'h106ed, 'h109be, 'h10bcd, 'h106fd, 'h1070d, 'h109bf, 'h1071d, 'h103bc, 'h1072d, 'h109c0, 'h1073d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074d, 'h109c1, 'h1075d, 'h1076d, 'h109c2, 'h1077d, 'h1078d, 'h109c3, 'h1079d, 'h10bcd, 'h107ad, 'h109c4, 'h107bd, 'h107cd, 'h109c5, 'h103bc, 'h107dd, 'h107ed, 'h109c6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fd, 'h1080d, 'h109c7, 'h1081d, 'h1082d, 'h109c8, 'h1083d, 'h1084d, 'h109c9, 'h10bcd, 'h1085d, 'h1086d, 'h109ca, 'h1087d, 'h103bc, 'h1088d, 'h109cb, 'h1089d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ad, 'h109cc, 'h108bd, 'h108cd, 'h109cd, 'h108dd, 'h106ed, 'h109ce, 'h10bdd, 'h106fd, 'h1070d, 'h109cf, 'h1071d, 'h1072d, 'h109d0, 'h103bc, 'h1073d, 'h1074d, 'h109d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075d, 'h1076d, 'h109d2, 'h1077d, 'h1078d, 'h109d3, 'h1079d, 'h10bdd, 'h107ad, 'h109d4, 'h107bd, 'h107cd, 'h109d5, 'h107dd, 'h103bc, 'h107ed, 'h109d6, 'h107fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080d, 'h109d7, 'h1081d, 'h1082d, 'h109d8, 'h1083d, 'h1084d, 'h109d9, 'h10bdd, 'h1085d, 'h1086d, 'h109da, 'h1087d, 'h1088d, 'h109db, 'h103bc, 'h1089d, 'h108ad, 'h109dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bd, 'h108cd, 'h109dd, 'h108dd, 'h106ed, 'h109de, 'h10bed, 'h106fd, 'h1070d, 'h109df, 'h1071d, 'h1072d, 'h109e0, 'h1073d, 'h103bc, 'h1074d, 'h109e1, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076d, 'h109e2, 'h1077d, 'h1078d, 'h109e3, 'h1079d, 'h10bed, 'h107ad, 'h109e4, 'h107bd, 'h107cd, 'h109e5, 'h107dd, 'h107ed, 'h109e6, 'h103bc, 'h107fd, 'h1080d, 'h109e7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081d, 'h1082d, 'h109e8, 'h1083d, 'h1084d, 'h109e9, 'h10bed, 'h1085d, 'h1086d, 'h109ea, 'h1087d, 'h1088d, 'h109eb, 'h1089d, 'h103bc, 'h108ad, 'h109ec, 'h108bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cd, 'h109ed, 'h108dd, 'h106ed, 'h109ee, 'h10bfd, 'h106fd, 'h1070d, 'h109ef, 'h1071d, 'h1072d, 'h109f0, 'h1073d, 'h1074d, 'h109f1, 'h103bc, 'h1075d, 'h1076d, 'h109f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077d, 'h1078d, 'h109f3, 'h1079d, 'h10bfd, 'h107ad, 'h109f4, 'h107bd, 'h107cd, 'h109f5, 'h107dd, 'h107ed, 'h109f6, 'h107fd, 'h103bc, 'h1080d, 'h109f7, 'h1081d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082d, 'h109f8, 'h1083d, 'h1084d, 'h109f9, 'h10bfd, 'h1085d, 'h1086d, 'h109fa, 'h1087d, 'h1088d, 'h109fb, 'h1089d, 'h108ad, 'h109fc, 'h103bc, 'h108bd, 'h108cd, 'h109fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dd, 'h106ed, 'h109fe, 'h10c0d, 'h106fd, 'h1070d, 'h109ff, 'h1071d, 'h1072d, 'h10a00, 'h1073d, 'h1074d, 'h10a01, 'h1075d, 'h103bc, 'h1076d, 'h10a02, 'h1077d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078d, 'h10a03, 'h1079d, 'h10c0d, 'h107ad, 'h10a04, 'h107bd, 'h107cd, 'h10a05, 'h107dd, 'h107ed, 'h10a06, 'h107fd, 'h1080d, 'h10a07, 'h103bc, 'h1081d, 'h1082d, 'h10a08, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083d, 'h1084d, 'h10a09, 'h10c0d, 'h1085d, 'h1086d, 'h10a0a, 'h1087d, 'h1088d, 'h10a0b, 'h1089d, 'h108ad, 'h10a0c, 'h108bd, 'h103bc, 'h108cd, 'h10a0d, 'h108dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ed, 'h10a0e, 'h10c1d, 'h106fd, 'h1070d, 'h10a0f, 'h1071d, 'h1072d, 'h10a10, 'h1073d, 'h1074d, 'h10a11, 'h1075d, 'h1076d, 'h10a12, 'h103bc, 'h1077d, 'h1078d, 'h10a13, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079d, 'h10c1d, 'h107ad, 'h10a14, 'h107bd, 'h107cd, 'h10a15, 'h107dd, 'h107ed, 'h10a16, 'h107fd, 'h1080d, 'h10a17, 'h1081d, 'h103bc, 'h1082d, 'h10a18, 'h1083d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084d, 'h10a19, 'h10c1d, 'h1085d, 'h1086d, 'h10a1a, 'h1087d, 'h1088d, 'h10a1b, 'h1089d, 'h108ad, 'h10a1c, 'h108bd, 'h108cd, 'h10a1d, 'h103bc, 'h108dd, 'h106ed, 'h10a1e, 'h10c2d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fd, 'h1070d, 'h10a1f, 'h1071d, 'h1072d, 'h10a20, 'h1073d, 'h1074d, 'h10a21, 'h1075d, 'h1076d, 'h10a22, 'h1077d, 'h103bc, 'h1078d, 'h10a23, 'h1079d, 'h10c2d, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ad, 'h10a24, 'h107bd, 'h107cd, 'h10a25, 'h107dd, 'h107ed, 'h10a26, 'h107fd, 'h1080d, 'h10a27, 'h1081d, 'h1082d, 'h10a28, 'h103bc, 'h1083d, 'h1084d, 'h10a29, 'h10c2d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085d, 'h1086d, 'h10a2a, 'h1087d, 'h1088d, 'h10a2b, 'h1089d, 'h108ad, 'h10a2c, 'h108bd, 'h108cd, 'h10a2d, 'h108dd, 'h103bc, 'h106ed, 'h10a2e, 'h10c3d, 'h106fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10a2f, 'h1071d, 'h1072d, 'h10a30, 'h1073d, 'h1074d, 'h10a31, 'h1075d, 'h1076d, 'h10a32, 'h1077d, 'h1078d, 'h10a33, 'h103bc, 'h1079d, 'h10c3d, 'h107ad, 'h10a34, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bd, 'h107cd, 'h10a35, 'h107dd, 'h107ed, 'h10a36, 'h107fd, 'h1080d, 'h10a37, 'h1081d, 'h1082d, 'h10a38, 'h1083d, 'h103bc, 'h1084d, 'h10a39, 'h10c3d, 'h1085d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086d, 'h10a3a, 'h1087d, 'h1088d, 'h10a3b, 'h1089d, 'h108ad, 'h10a3c, 'h108bd, 'h108cd, 'h10a3d, 'h108dd, 'h106ed, 'h10a3e, 'h10c4d, 'h103bc, 'h106fd, 'h1070d, 'h10a3f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071d, 'h1072d, 'h10a40, 'h1073d, 'h1074d, 'h10a41, 'h1075d, 'h1076d, 'h10a42, 'h1077d, 'h1078d, 'h10a43, 'h1079d, 'h10c4d, 'h103bc, 'h107ad, 'h10a44, 'h107bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cd, 'h10a45, 'h107dd, 'h107ed, 'h10a46, 'h107fd, 'h1080d, 'h10a47, 'h1081d, 'h1082d, 'h10a48, 'h1083d, 'h1084d, 'h10a49, 'h10c4d, 'h103bc, 'h1085d, 'h1086d, 'h10a4a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087d, 'h1088d, 'h10a4b, 'h1089d, 'h108ad, 'h10a4c, 'h108bd, 'h108cd, 'h10a4d, 'h108dd, 'h106ed, 'h10a4e, 'h10c5d, 'h106fd, 'h103bc, 'h1070d, 'h10a4f, 'h1071d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072d, 'h10a50, 'h1073d, 'h1074d, 'h10a51, 'h1075d, 'h1076d, 'h10a52, 'h1077d, 'h1078d, 'h10a53, 'h1079d, 'h10c5d, 'h107ad, 'h10a54, 'h103bc, 'h107bd, 'h107cd, 'h10a55, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dd, 'h107ed, 'h10a56, 'h107fd, 'h1080d, 'h10a57, 'h1081d, 'h1082d, 'h10a58, 'h1083d, 'h1084d, 'h10a59, 'h10c5d, 'h1085d, 'h103bc, 'h1086d, 'h10a5a, 'h1087d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088d, 'h10a5b, 'h1089d, 'h108ad, 'h10a5c, 'h108bd, 'h108cd, 'h10a5d, 'h108dd, 'h106ed, 'h10a5e, 'h10c6d, 'h106fd, 'h1070d, 'h10a5f, 'h103bc, 'h1071d, 'h1072d, 'h10a60, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h1074d, 'h10a61, 'h1075d, 'h1076d, 'h10a62, 'h1077d, 'h1078d, 'h10a63, 'h1079d, 'h10c6d, 'h107ad, 'h10a64, 'h107bd, 'h103bc, 'h107cd, 'h10a65, 'h107dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ed, 'h10a66, 'h107fd, 'h1080d, 'h10a67, 'h1081d, 'h1082d, 'h10a68, 'h1083d, 'h1084d, 'h10a69, 'h10c6d, 'h1085d, 'h1086d, 'h10a6a, 'h103bc, 'h1087d, 'h1088d, 'h10a6b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089d, 'h108ad, 'h10a6c, 'h108bd, 'h108cd, 'h10a6d, 'h108dd, 'h106ed, 'h10a6e, 'h10c7d, 'h106fd, 'h1070d, 'h10a6f, 'h1071d, 'h103bc, 'h1072d, 'h10a70, 'h1073d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074d, 'h10a71, 'h1075d, 'h1076d, 'h10a72, 'h1077d, 'h1078d, 'h10a73, 'h1079d, 'h10c7d, 'h107ad, 'h10a74, 'h107bd, 'h107cd, 'h10a75, 'h103bc, 'h107dd, 'h107ed, 'h10a76, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fd, 'h1080d, 'h10a77, 'h1081d, 'h1082d, 'h10a78, 'h1083d, 'h1084d, 'h10a79, 'h10c7d, 'h1085d, 'h1086d, 'h10a7a, 'h1087d, 'h103bc, 'h1088d, 'h10a7b, 'h1089d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ad, 'h10a7c, 'h108bd, 'h108cd, 'h10a7d, 'h108dd, 'h106ed, 'h10a7e, 'h10c8d, 'h106fd, 'h1070d, 'h10a7f, 'h1071d, 'h1072d, 'h10a80, 'h103bc, 'h1073d, 'h1074d, 'h10a81, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075d, 'h1076d, 'h10a82, 'h1077d, 'h1078d, 'h10a83, 'h1079d, 'h10c8d, 'h107ad, 'h10a84, 'h107bd, 'h107cd, 'h10a85, 'h107dd, 'h103bc, 'h107ed, 'h10a86, 'h107fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080d, 'h10a87, 'h1081d, 'h1082d, 'h10a88, 'h1083d, 'h1084d, 'h10a89, 'h10c8d, 'h1085d, 'h1086d, 'h10a8a, 'h1087d, 'h1088d, 'h10a8b, 'h103bc, 'h1089d, 'h108ad, 'h10a8c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bd, 'h108cd, 'h10a8d, 'h108dd, 'h106ed, 'h10a8e, 'h10c9d, 'h106fd, 'h1070d, 'h10a8f, 'h1071d, 'h1072d, 'h10a90, 'h1073d, 'h103bc, 'h1074d, 'h10a91, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076d, 'h10a92, 'h1077d, 'h1078d, 'h10a93, 'h1079d, 'h10c9d, 'h107ad, 'h10a94, 'h107bd, 'h107cd, 'h10a95, 'h107dd, 'h107ed, 'h10a96, 'h103bc, 'h107fd, 'h1080d, 'h10a97, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081d, 'h1082d, 'h10a98, 'h1083d, 'h1084d, 'h10a99, 'h10c9d, 'h1085d, 'h1086d, 'h10a9a, 'h1087d, 'h1088d, 'h10a9b, 'h1089d, 'h103bc, 'h108ad, 'h10a9c, 'h108bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cd, 'h10a9d, 'h108dd, 'h106ed, 'h10a9e, 'h10cad, 'h106fd, 'h1070d, 'h10a9f, 'h1071d, 'h1072d, 'h10aa0, 'h1073d, 'h1074d, 'h10aa1, 'h103bc, 'h1075d, 'h1076d, 'h10aa2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077d, 'h1078d, 'h10aa3, 'h1079d, 'h10cad, 'h107ad, 'h10aa4, 'h107bd, 'h107cd, 'h10aa5, 'h107dd, 'h107ed, 'h10aa6, 'h107fd, 'h103bc, 'h1080d, 'h10aa7, 'h1081d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082d, 'h10aa8, 'h1083d, 'h1084d, 'h10aa9, 'h10cad, 'h1085d, 'h1086d, 'h10aaa, 'h1087d, 'h1088d, 'h10aab, 'h1089d, 'h108ad, 'h10aac, 'h103bc, 'h108bd, 'h108cd, 'h10aad, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dd, 'h106ed, 'h10aae, 'h10cbd, 'h106fd, 'h1070d, 'h10aaf, 'h1071d, 'h1072d, 'h10ab0, 'h1073d, 'h1074d, 'h10ab1, 'h1075d, 'h103bc, 'h1076d, 'h10ab2, 'h1077d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078d, 'h10ab3, 'h1079d, 'h10cbd, 'h107ad, 'h10ab4, 'h107bd, 'h107cd, 'h10ab5, 'h107dd, 'h107ed, 'h10ab6, 'h107fd, 'h1080d, 'h10ab7, 'h103bc, 'h1081d, 'h1082d, 'h10ab8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083d, 'h1084d, 'h10ab9, 'h10cbd, 'h1085d, 'h1086d, 'h10aba, 'h1087d, 'h1088d, 'h10abb, 'h1089d, 'h108ad, 'h10abc, 'h108bd, 'h103bc, 'h108cd, 'h10abd, 'h108dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ed, 'h10abe, 'h10ccd, 'h106fd, 'h1070d, 'h10abf, 'h1071d, 'h1072d, 'h10ac0, 'h1073d, 'h1074d, 'h10ac1, 'h1075d, 'h1076d, 'h10ac2, 'h103bc, 'h1077d, 'h1078d, 'h10ac3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079d, 'h10ccd, 'h107ad, 'h10ac4, 'h107bd, 'h107cd, 'h10ac5, 'h107dd, 'h107ed, 'h10ac6, 'h107fd, 'h1080d, 'h10ac7, 'h1081d, 'h103bc, 'h1082d, 'h10ac8, 'h1083d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084d, 'h10ac9, 'h10ccd, 'h1085d, 'h1086d, 'h10aca, 'h1087d, 'h1088d, 'h10acb, 'h1089d, 'h108ad, 'h10acc, 'h108bd, 'h108cd, 'h10acd, 'h103bc, 'h108dd, 'h106ed, 'h10ace, 'h10cdd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fd, 'h1070d, 'h10acf, 'h1071d, 'h1072d, 'h10ad0, 'h1073d, 'h1074d, 'h10ad1, 'h1075d, 'h1076d, 'h10ad2, 'h1077d, 'h103bc, 'h1078d, 'h10ad3, 'h1079d, 'h10cdd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ad, 'h10ad4, 'h107bd, 'h107cd, 'h10ad5, 'h107dd, 'h107ed, 'h10ad6, 'h107fd, 'h1080d, 'h10ad7, 'h1081d, 'h1082d, 'h10ad8, 'h103bc, 'h1083d, 'h1084d, 'h10ad9, 'h10cdd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085d, 'h1086d, 'h10ada, 'h1087d, 'h1088d, 'h10adb, 'h1089d, 'h108ad, 'h10adc, 'h108bd, 'h108cd, 'h10add, 'h108dd, 'h103bc, 'h106ed, 'h108de, 'h10aed, 'h106fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h108df, 'h1071d, 'h1072d, 'h108e0, 'h1073d, 'h1074d, 'h108e1, 'h1075d, 'h1076d, 'h108e2, 'h1077d, 'h1078d, 'h108e3, 'h103bc, 'h1079d, 'h10aed, 'h107ad, 'h108e4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bd, 'h107cd, 'h108e5, 'h107dd, 'h107ed, 'h108e6, 'h107fd, 'h1080d, 'h108e7, 'h1081d, 'h1082d, 'h108e8, 'h1083d, 'h103bc, 'h1084d, 'h108e9, 'h10aed, 'h1085d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086d, 'h108ea, 'h1087d, 'h1088d, 'h108eb, 'h1089d, 'h108ad, 'h108ec, 'h108bd, 'h108cd, 'h108ed, 'h108dd, 'h106ed, 'h108ee, 'h10afd, 'h103bc, 'h106fd, 'h1070d, 'h108ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071d, 'h1072d, 'h108f0, 'h1073d, 'h1074d, 'h108f1, 'h1075d, 'h1076d, 'h108f2, 'h1077d, 'h1078d, 'h108f3, 'h1079d, 'h10afd, 'h103bc, 'h107ad, 'h108f4, 'h107bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cd, 'h108f5, 'h107dd, 'h107ed, 'h108f6, 'h107fd, 'h1080d, 'h108f7, 'h1081d, 'h1082d, 'h108f8, 'h1083d, 'h1084d, 'h108f9, 'h10afd, 'h103bc, 'h1085d, 'h1086d, 'h108fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087d, 'h1088d, 'h108fb, 'h1089d, 'h108ad, 'h108fc, 'h108bd, 'h108cd, 'h108fd, 'h108dd, 'h106ed, 'h108fe, 'h10b0d, 'h106fd, 'h103bc, 'h1070d, 'h108ff, 'h1071d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072d, 'h10900, 'h1073d, 'h1074d, 'h10901, 'h1075d, 'h1076d, 'h10902, 'h1077d, 'h1078d, 'h10903, 'h1079d, 'h10b0d, 'h107ad, 'h10904, 'h103bc, 'h107bd, 'h107cd, 'h10905, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dd, 'h107ed, 'h10906, 'h107fd, 'h1080d, 'h10907, 'h1081d, 'h1082d, 'h10908, 'h1083d, 'h1084d, 'h10909, 'h10b0d, 'h1085d, 'h103bc, 'h1086d, 'h1090a, 'h1087d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088d, 'h1090b, 'h1089d, 'h108ad, 'h1090c, 'h108bd, 'h108cd, 'h1090d, 'h108dd, 'h106ed, 'h1090e, 'h10b1d, 'h106fd, 'h1070d, 'h1090f, 'h103bc, 'h1071d, 'h1072d, 'h10910, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h1074d, 'h10911, 'h1075d, 'h1076d, 'h10912, 'h1077d, 'h1078d, 'h10913, 'h1079d, 'h10b1d, 'h107ad, 'h10914, 'h107bd, 'h103bc, 'h107cd, 'h10915, 'h107dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ed, 'h10916, 'h107fd, 'h1080d, 'h10917, 'h1081d, 'h1082d, 'h10918, 'h1083d, 'h1084d, 'h10919, 'h10b1d, 'h1085d, 'h1086d, 'h1091a, 'h103bc, 'h1087d, 'h1088d, 'h1091b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089d, 'h108ad, 'h1091c, 'h108bd, 'h108cd, 'h1091d, 'h108dd, 'h106ed, 'h1091e, 'h10b2d, 'h106fd, 'h1070d, 'h1091f, 'h1071d, 'h103bc, 'h1072d, 'h10920, 'h1073d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074d, 'h10921, 'h1075d, 'h1076d, 'h10922, 'h1077d, 'h1078d, 'h10923, 'h1079d, 'h10b2d, 'h107ad, 'h10924, 'h107bd, 'h107cd, 'h10925, 'h103bc, 'h107dd, 'h107ed, 'h10926, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fd, 'h1080d, 'h10927, 'h1081d, 'h1082d, 'h10928, 'h1083d, 'h1084d, 'h10929, 'h10b2d, 'h1085d, 'h1086d, 'h1092a, 'h1087d, 'h103bc, 'h1088d, 'h1092b, 'h1089d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ad, 'h1092c, 'h108bd, 'h108cd, 'h1092d, 'h108dd, 'h106ed, 'h1092e, 'h10b3d, 'h106fd, 'h1070d, 'h1092f, 'h1071d, 'h1072d, 'h10930, 'h103bc, 'h1073d, 'h1074d, 'h10931, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075d, 'h1076d, 'h10932, 'h1077d, 'h1078d, 'h10933, 'h1079d, 'h10b3d, 'h107ad, 'h10934, 'h107bd, 'h107cd, 'h10935, 'h107dd, 'h103bc, 'h107ed, 'h10936, 'h107fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080d, 'h10937, 'h1081d, 'h1082d, 'h10938, 'h1083d, 'h1084d, 'h10939, 'h10b3d, 'h1085d, 'h1086d, 'h1093a, 'h1087d, 'h1088d, 'h1093b, 'h103bc, 'h1089d, 'h108ad, 'h1093c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bd, 'h108cd, 'h1093d, 'h108dd, 'h106ed, 'h1093e, 'h10b4d, 'h106fd, 'h1070d, 'h1093f, 'h1071d, 'h1072d, 'h10940, 'h1073d, 'h103bc, 'h1074d, 'h10941, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076d, 'h10942, 'h1077d, 'h1078d, 'h10943, 'h1079d, 'h10b4d, 'h107ad, 'h10944, 'h107bd, 'h107cd, 'h10945, 'h107dd, 'h107ed, 'h10946, 'h103bc, 'h107fd, 'h1080d, 'h10947, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081d, 'h1082d, 'h10948, 'h1083d, 'h1084d, 'h10949, 'h10b4d, 'h1085d, 'h1086d, 'h1094a, 'h1087d, 'h1088d, 'h1094b, 'h1089d, 'h103bc, 'h108ad, 'h1094c, 'h108bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cd, 'h1094d, 'h108dd, 'h106ed, 'h1094e, 'h10b5d, 'h106fd, 'h1070d, 'h1094f, 'h1071d, 'h1072d, 'h10950, 'h1073d, 'h1074d, 'h10951, 'h103bc, 'h1075d, 'h1076d, 'h10952, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077d, 'h1078d, 'h10953, 'h1079d, 'h10b5d, 'h107ad, 'h10954, 'h107bd, 'h107cd, 'h10955, 'h107dd, 'h107ed, 'h10956, 'h107fd, 'h103bc, 'h1080d, 'h10957, 'h1081d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082d, 'h10958, 'h1083d, 'h1084d, 'h10959, 'h10b5d, 'h1085d, 'h1086d, 'h1095a, 'h1087d, 'h1088d, 'h1095b, 'h1089d, 'h108ad, 'h1095c, 'h103bc, 'h108bd, 'h108cd, 'h1095d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dd, 'h106ed, 'h1095e, 'h10b6d, 'h106fd, 'h1070d, 'h1095f, 'h1071d, 'h1072d, 'h10960, 'h1073d, 'h1074d, 'h10961, 'h1075d, 'h103bc, 'h1076d, 'h10962, 'h1077d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078d, 'h10963, 'h1079d, 'h10b6d, 'h107ad, 'h10964, 'h107bd, 'h107cd, 'h10965, 'h107dd, 'h107ed, 'h10966, 'h107fd, 'h1080d, 'h10967, 'h103bc, 'h1081d, 'h1082d, 'h10968, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083d, 'h1084d, 'h10969, 'h10b6d, 'h1085d, 'h1086d, 'h1096a, 'h1087d, 'h1088d, 'h1096b, 'h1089d, 'h108ad, 'h1096c, 'h108bd, 'h103bc, 'h108cd, 'h1096d, 'h108dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ed, 'h1096e, 'h10b7d, 'h106fd, 'h1070d, 'h1096f, 'h1071d, 'h1072d, 'h10970, 'h1073d, 'h1074d, 'h10971, 'h1075d, 'h1076d, 'h10972, 'h103bc, 'h1077d, 'h1078d, 'h10973, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079d, 'h10b7d, 'h107ad, 'h10974, 'h107bd, 'h107cd, 'h10975, 'h107dd, 'h107ed, 'h10976, 'h107fd, 'h1080d, 'h10977, 'h1081d, 'h103bc, 'h1082d, 'h10978, 'h1083d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084d, 'h10979, 'h10b7d, 'h1085d, 'h1086d, 'h1097a, 'h1087d, 'h1088d, 'h1097b, 'h1089d, 'h108ad, 'h1097c, 'h108bd, 'h108cd, 'h1097d, 'h103bc, 'h108dd, 'h106ed, 'h1097e, 'h10b8d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fd, 'h1070d, 'h1097f, 'h1071d, 'h1072d, 'h10980, 'h1073d, 'h1074d, 'h10981, 'h1075d, 'h1076d, 'h10982, 'h1077d, 'h103bc, 'h1078d, 'h10983, 'h1079d, 'h10b8d, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ad, 'h10984, 'h107bd, 'h107cd, 'h10985, 'h107dd, 'h107ed, 'h10986, 'h107fd, 'h1080d, 'h10987, 'h1081d, 'h1082d, 'h10988, 'h103bc, 'h1083d, 'h1084d, 'h10989, 'h10b8d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085d, 'h1086d, 'h1098a, 'h1087d, 'h1088d, 'h1098b, 'h1089d, 'h108ad, 'h1098c, 'h108bd, 'h108cd, 'h1098d, 'h108dd, 'h103bc, 'h106ed, 'h1098e, 'h10b9d, 'h106fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h1098f, 'h1071d, 'h1072d, 'h10990, 'h1073d, 'h1074d, 'h10991, 'h1075d, 'h1076d, 'h10992, 'h1077d, 'h1078d, 'h10993, 'h103bc, 'h1079d, 'h10b9d, 'h107ad, 'h10994, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bd, 'h107cd, 'h10995, 'h107dd, 'h107ed, 'h10996, 'h107fd, 'h1080d, 'h10997, 'h1081d, 'h1082d, 'h10998, 'h1083d, 'h103bc, 'h1084d, 'h10999, 'h10b9d, 'h1085d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086d, 'h1099a, 'h1087d, 'h1088d, 'h1099b, 'h1089d, 'h108ad, 'h1099c, 'h108bd, 'h108cd, 'h1099d, 'h108dd, 'h106ed, 'h1099e, 'h10bad, 'h103bc, 'h106fd, 'h1070d, 'h1099f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071d, 'h1072d, 'h109a0, 'h1073d, 'h1074d, 'h109a1, 'h1075d, 'h1076d, 'h109a2, 'h1077d, 'h1078d, 'h109a3, 'h1079d, 'h10bad, 'h103bc, 'h107ad, 'h109a4, 'h107bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cd, 'h109a5, 'h107dd, 'h107ed, 'h109a6, 'h107fd, 'h1080d, 'h109a7, 'h1081d, 'h1082d, 'h109a8, 'h1083d, 'h1084d, 'h109a9, 'h10bad, 'h103bc, 'h1085d, 'h1086d, 'h109aa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087d, 'h1088d, 'h109ab, 'h1089d, 'h108ad, 'h109ac, 'h108bd, 'h108cd, 'h109ad, 'h108dd, 'h106ed, 'h109ae, 'h10bbd, 'h106fd, 'h103bc, 'h1070d, 'h109af, 'h1071d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072d, 'h109b0, 'h1073d, 'h1074d, 'h109b1, 'h1075d, 'h1076d, 'h109b2, 'h1077d, 'h1078d, 'h109b3, 'h1079d, 'h10bbd, 'h107ad, 'h109b4, 'h103bc, 'h107bd, 'h107cd, 'h109b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dd, 'h107ed, 'h109b6, 'h107fd, 'h1080d, 'h109b7, 'h1081d, 'h1082d, 'h109b8, 'h1083d, 'h1084d, 'h109b9, 'h10bbd, 'h1085d, 'h103bc, 'h1086d, 'h109ba, 'h1087d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088d, 'h109bb, 'h1089d, 'h108ad, 'h109bc, 'h108bd, 'h108cd, 'h109bd, 'h108dd, 'h106ed, 'h109be, 'h10bcd, 'h106fd, 'h1070d, 'h109bf, 'h103bc, 'h1071d, 'h1072d, 'h109c0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h1074d, 'h109c1, 'h1075d, 'h1076d, 'h109c2, 'h1077d, 'h1078d, 'h109c3, 'h1079d, 'h10bcd, 'h107ad, 'h109c4, 'h107bd, 'h103bc, 'h107cd, 'h109c5, 'h107dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ed, 'h109c6, 'h107fd, 'h1080d, 'h109c7, 'h1081d, 'h1082d, 'h109c8, 'h1083d, 'h1084d, 'h109c9, 'h10bcd, 'h1085d, 'h1086d, 'h109ca, 'h103bc, 'h1087d, 'h1088d, 'h109cb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089d, 'h108ad, 'h109cc, 'h108bd, 'h108cd, 'h109cd, 'h108dd, 'h106ed, 'h109ce, 'h10bdd, 'h106fd, 'h1070d, 'h109cf, 'h1071d, 'h103bc, 'h1072d, 'h109d0, 'h1073d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074d, 'h109d1, 'h1075d, 'h1076d, 'h109d2, 'h1077d, 'h1078d, 'h109d3, 'h1079d, 'h10bdd, 'h107ad, 'h109d4, 'h107bd, 'h107cd, 'h109d5, 'h103bc, 'h107dd, 'h107ed, 'h109d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fd, 'h1080d, 'h109d7, 'h1081d, 'h1082d, 'h109d8, 'h1083d, 'h1084d, 'h109d9, 'h10bdd, 'h1085d, 'h1086d, 'h109da, 'h1087d, 'h103bc, 'h1088d, 'h109db, 'h1089d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ad, 'h109dc, 'h108bd, 'h108cd, 'h109dd, 'h108dd, 'h106ed, 'h109de, 'h10bed, 'h106fd, 'h1070d, 'h109df, 'h1071d, 'h1072d, 'h109e0, 'h103bc, 'h1073d, 'h1074d, 'h109e1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075d, 'h1076d, 'h109e2, 'h1077d, 'h1078d, 'h109e3, 'h1079d, 'h10bed, 'h107ad, 'h109e4, 'h107bd, 'h107cd, 'h109e5, 'h107dd, 'h103bc, 'h107ed, 'h109e6, 'h107fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080d, 'h109e7, 'h1081d, 'h1082d, 'h109e8, 'h1083d, 'h1084d, 'h109e9, 'h10bed, 'h1085d, 'h1086d, 'h109ea, 'h1087d, 'h1088d, 'h109eb, 'h103bc, 'h1089d, 'h108ad, 'h109ec, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bd, 'h108cd, 'h109ed, 'h108dd, 'h106ed, 'h109ee, 'h10bfd, 'h106fd, 'h1070d, 'h109ef, 'h1071d, 'h1072d, 'h109f0, 'h1073d, 'h103bc, 'h1074d, 'h109f1, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076d, 'h109f2, 'h1077d, 'h1078d, 'h109f3, 'h1079d, 'h10bfd, 'h107ad, 'h109f4, 'h107bd, 'h107cd, 'h109f5, 'h107dd, 'h107ed, 'h109f6, 'h103bc, 'h107fd, 'h1080d, 'h109f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081d, 'h1082d, 'h109f8, 'h1083d, 'h1084d, 'h109f9, 'h10bfd, 'h1085d, 'h1086d, 'h109fa, 'h1087d, 'h1088d, 'h109fb, 'h1089d, 'h103bc, 'h108ad, 'h109fc, 'h108bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cd, 'h109fd, 'h108dd, 'h106ed, 'h109fe, 'h10c0d, 'h106fd, 'h1070d, 'h109ff, 'h1071d, 'h1072d, 'h10a00, 'h1073d, 'h1074d, 'h10a01, 'h103bc, 'h1075d, 'h1076d, 'h10a02, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077d, 'h1078d, 'h10a03, 'h1079d, 'h10c0d, 'h107ad, 'h10a04, 'h107bd, 'h107cd, 'h10a05, 'h107dd, 'h107ed, 'h10a06, 'h107fd, 'h103bc, 'h1080d, 'h10a07, 'h1081d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082d, 'h10a08, 'h1083d, 'h1084d, 'h10a09, 'h10c0d, 'h1085d, 'h1086d, 'h10a0a, 'h1087d, 'h1088d, 'h10a0b, 'h1089d, 'h108ad, 'h10a0c, 'h103bc, 'h108bd, 'h108cd, 'h10a0d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dd, 'h106ed, 'h10a0e, 'h10c1d, 'h106fd, 'h1070d, 'h10a0f, 'h1071d, 'h1072d, 'h10a10, 'h1073d, 'h1074d, 'h10a11, 'h1075d, 'h103bc, 'h1076d, 'h10a12, 'h1077d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078d, 'h10a13, 'h1079d, 'h10c1d, 'h107ad, 'h10a14, 'h107bd, 'h107cd, 'h10a15, 'h107dd, 'h107ed, 'h10a16, 'h107fd, 'h1080d, 'h10a17, 'h103bc, 'h1081d, 'h1082d, 'h10a18, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083d, 'h1084d, 'h10a19, 'h10c1d, 'h1085d, 'h1086d, 'h10a1a, 'h1087d, 'h1088d, 'h10a1b, 'h1089d, 'h108ad, 'h10a1c, 'h108bd, 'h103bc, 'h108cd, 'h10a1d, 'h108dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ed, 'h10a1e, 'h10c2d, 'h106fd, 'h1070d, 'h10a1f, 'h1071d, 'h1072d, 'h10a20, 'h1073d, 'h1074d, 'h10a21, 'h1075d, 'h1076d, 'h10a22, 'h103bc, 'h1077d, 'h1078d, 'h10a23, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079d, 'h10c2d, 'h107ad, 'h10a24, 'h107bd, 'h107cd, 'h10a25, 'h107dd, 'h107ed, 'h10a26, 'h107fd, 'h1080d, 'h10a27, 'h1081d, 'h103bc, 'h1082d, 'h10a28, 'h1083d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084d, 'h10a29, 'h10c2d, 'h1085d, 'h1086d, 'h10a2a, 'h1087d, 'h1088d, 'h10a2b, 'h1089d, 'h108ad, 'h10a2c, 'h108bd, 'h108cd, 'h10a2d, 'h103bc, 'h108dd, 'h106ed, 'h10a2e, 'h10c3d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fd, 'h1070d, 'h10a2f, 'h1071d, 'h1072d, 'h10a30, 'h1073d, 'h1074d, 'h10a31, 'h1075d, 'h1076d, 'h10a32, 'h1077d, 'h103bc, 'h1078d, 'h10a33, 'h1079d, 'h10c3d, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ad, 'h10a34, 'h107bd, 'h107cd, 'h10a35, 'h107dd, 'h107ed, 'h10a36, 'h107fd, 'h1080d, 'h10a37, 'h1081d, 'h1082d, 'h10a38, 'h103bc, 'h1083d, 'h1084d, 'h10a39, 'h10c3d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085d, 'h1086d, 'h10a3a, 'h1087d, 'h1088d, 'h10a3b, 'h1089d, 'h108ad, 'h10a3c, 'h108bd, 'h108cd, 'h10a3d, 'h108dd, 'h103bc, 'h106ed, 'h10a3e, 'h10c4d, 'h106fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10a3f, 'h1071d, 'h1072d, 'h10a40, 'h1073d, 'h1074d, 'h10a41, 'h1075d, 'h1076d, 'h10a42, 'h1077d, 'h1078d, 'h10a43, 'h103bc, 'h1079d, 'h10c4d, 'h107ad, 'h10a44, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bd, 'h107cd, 'h10a45, 'h107dd, 'h107ed, 'h10a46, 'h107fd, 'h1080d, 'h10a47, 'h1081d, 'h1082d, 'h10a48, 'h1083d, 'h103bc, 'h1084d, 'h10a49, 'h10c4d, 'h1085d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086d, 'h10a4a, 'h1087d, 'h1088d, 'h10a4b, 'h1089d, 'h108ad, 'h10a4c, 'h108bd, 'h108cd, 'h10a4d, 'h108dd, 'h106ed, 'h10a4e, 'h10c5d, 'h103bc, 'h106fd, 'h1070d, 'h10a4f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071d, 'h1072d, 'h10a50, 'h1073d, 'h1074d, 'h10a51, 'h1075d, 'h1076d, 'h10a52, 'h1077d, 'h1078d, 'h10a53, 'h1079d, 'h10c5d, 'h103bc, 'h107ad, 'h10a54, 'h107bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cd, 'h10a55, 'h107dd, 'h107ed, 'h10a56, 'h107fd, 'h1080d, 'h10a57, 'h1081d, 'h1082d, 'h10a58, 'h1083d, 'h1084d, 'h10a59, 'h10c5d, 'h103bc, 'h1085d, 'h1086d, 'h10a5a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087d, 'h1088d, 'h10a5b, 'h1089d, 'h108ad, 'h10a5c, 'h108bd, 'h108cd, 'h10a5d, 'h108dd, 'h106ed, 'h10a5e, 'h10c6d, 'h106fd, 'h103bc, 'h1070d, 'h10a5f, 'h1071d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072d, 'h10a60, 'h1073d, 'h1074d, 'h10a61, 'h1075d, 'h1076d, 'h10a62, 'h1077d, 'h1078d, 'h10a63, 'h1079d, 'h10c6d, 'h107ad, 'h10a64, 'h103bc, 'h107bd, 'h107cd, 'h10a65, 'h21f8e, 'h21f8f, 'h21f8d, 'h107dd, 'h107ed, 'h10a66, 'h107fd, 'h1080d, 'h10a67, 'h1081d, 'h1082d, 'h10a68, 'h1083d, 'h1084d, 'h10a69, 'h10c6d, 'h1085d, 'h103bc, 'h1086d, 'h10a6a, 'h1087d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088d, 'h10a6b, 'h1089d, 'h108ad, 'h10a6c, 'h108bd, 'h108cd, 'h10a6d, 'h108dd, 'h106ed, 'h10a6e, 'h10c7d, 'h106fd, 'h1070d, 'h10a6f, 'h103bc, 'h1071d, 'h1072d, 'h10a70, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h1074d, 'h10a71, 'h1075d, 'h1076d, 'h10a72, 'h1077d, 'h1078d, 'h10a73, 'h1079d, 'h10c7d, 'h107ad, 'h10a74, 'h107bd, 'h103bc, 'h107cd, 'h10a75, 'h107dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ed, 'h10a76, 'h107fd, 'h1080d, 'h10a77, 'h1081d, 'h1082d, 'h10a78, 'h1083d, 'h1084d, 'h10a79, 'h10c7d, 'h1085d, 'h1086d, 'h10a7a, 'h103bc, 'h1087d, 'h1088d, 'h10a7b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089d, 'h108ad, 'h10a7c, 'h108bd, 'h108cd, 'h10a7d, 'h108dd, 'h106ed, 'h10a7e, 'h10c8d, 'h106fd, 'h1070d, 'h10a7f, 'h1071d, 'h103bc, 'h1072d, 'h10a80, 'h1073d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074d, 'h10a81, 'h1075d, 'h1076d, 'h10a82, 'h1077d, 'h1078d, 'h10a83, 'h1079d, 'h10c8d, 'h107ad, 'h10a84, 'h107bd, 'h107cd, 'h10a85, 'h103bc, 'h107dd, 'h107ed, 'h10a86, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fd, 'h1080d, 'h10a87, 'h1081d, 'h1082d, 'h10a88, 'h1083d, 'h1084d, 'h10a89, 'h10c8d, 'h1085d, 'h1086d, 'h10a8a, 'h1087d, 'h103bc, 'h1088d, 'h10a8b, 'h1089d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ad, 'h10a8c, 'h108bd, 'h108cd, 'h10a8d, 'h108dd, 'h106ed, 'h10a8e, 'h10c9d, 'h106fd, 'h1070d, 'h10a8f, 'h1071d, 'h1072d, 'h10a90, 'h103bc, 'h1073d, 'h1074d, 'h10a91, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075d, 'h1076d, 'h10a92, 'h1077d, 'h1078d, 'h10a93, 'h1079d, 'h10c9d, 'h107ad, 'h10a94, 'h107bd, 'h107cd, 'h10a95, 'h107dd, 'h103bc, 'h107ed, 'h10a96, 'h107fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080d, 'h10a97, 'h1081d, 'h1082d, 'h10a98, 'h1083d, 'h1084d, 'h10a99, 'h10c9d, 'h1085d, 'h1086d, 'h10a9a, 'h1087d, 'h1088d, 'h10a9b, 'h103bc, 'h1089d, 'h108ad, 'h10a9c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bd, 'h108cd, 'h10a9d, 'h108dd, 'h106ed, 'h10a9e, 'h10cad, 'h106fd, 'h1070d, 'h10a9f, 'h1071d, 'h1072d, 'h10aa0, 'h1073d, 'h103bc, 'h1074d, 'h10aa1, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076d, 'h10aa2, 'h1077d, 'h1078d, 'h10aa3, 'h1079d, 'h10cad, 'h107ad, 'h10aa4, 'h107bd, 'h107cd, 'h10aa5, 'h107dd, 'h107ed, 'h10aa6, 'h103bc, 'h107fd, 'h1080d, 'h10aa7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081d, 'h1082d, 'h10aa8, 'h1083d, 'h1084d, 'h10aa9, 'h10cad, 'h1085d, 'h1086d, 'h10aaa, 'h1087d, 'h1088d, 'h10aab, 'h1089d, 'h103bc, 'h108ad, 'h10aac, 'h108bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cd, 'h10aad, 'h108dd, 'h106ed, 'h10aae, 'h10cbd, 'h106fd, 'h1070d, 'h10aaf, 'h1071d, 'h1072d, 'h10ab0, 'h1073d, 'h1074d, 'h10ab1, 'h103bc, 'h1075d, 'h1076d, 'h10ab2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077d, 'h1078d, 'h10ab3, 'h1079d, 'h10cbd, 'h107ad, 'h10ab4, 'h107bd, 'h107cd, 'h10ab5, 'h107dd, 'h107ed, 'h10ab6, 'h107fd, 'h103bc, 'h1080d, 'h10ab7, 'h1081d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082d, 'h10ab8, 'h1083d, 'h1084d, 'h10ab9, 'h10cbd, 'h1085d, 'h1086d, 'h10aba, 'h1087d, 'h1088d, 'h10abb, 'h1089d, 'h108ad, 'h10abc, 'h103bc, 'h108bd, 'h108cd, 'h10abd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dd, 'h106ed, 'h10abe, 'h10ccd, 'h106fd, 'h1070d, 'h10abf, 'h1071d, 'h1072d, 'h10ac0, 'h1073d, 'h1074d, 'h10ac1, 'h1075d, 'h103bc, 'h1076d, 'h10ac2, 'h1077d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078d, 'h10ac3, 'h1079d, 'h10ccd, 'h107ad, 'h10ac4, 'h107bd, 'h107cd, 'h10ac5, 'h107dd, 'h107ed, 'h10ac6, 'h107fd, 'h1080d, 'h10ac7, 'h103bc, 'h1081d, 'h1082d, 'h10ac8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083d, 'h1084d, 'h10ac9, 'h10ccd, 'h1085d, 'h1086d, 'h10aca, 'h1087d, 'h1088d, 'h10acb, 'h1089d, 'h108ad, 'h10acc, 'h108bd, 'h103bc, 'h108cd, 'h10acd, 'h108dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ed, 'h10ace, 'h10cdd, 'h106fd, 'h1070d, 'h10acf, 'h1071d, 'h1072d, 'h10ad0, 'h1073d, 'h1074d, 'h10ad1, 'h1075d, 'h1076d, 'h10ad2, 'h103bc, 'h1077d, 'h1078d, 'h10ad3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079d, 'h10cdd, 'h107ad, 'h10ad4, 'h107bd, 'h107cd, 'h10ad5, 'h107dd, 'h107ed, 'h10ad6, 'h107fd, 'h1080d, 'h10ad7, 'h1081d, 'h103bc, 'h1082d, 'h10ad8, 'h1083d, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084d, 'h10ad9, 'h10cdd, 'h1085d, 'h1086d, 'h10ada, 'h1087d, 'h1088d, 'h10adb, 'h1089d, 'h108ad, 'h10adc, 'h108bd, 'h108cd, 'h10add, 'h103bc, 'h108dd, 'h21f8c, 'h21f8b, 'h21f8f, 'h10440, 'h21f8d, 'h21f8a, 'h10443, 'h10442, 'h1043f, 'h10441, 'h103dc, 'h103dd, 'h21f88, 'h21f89, 'h21f87, 'h103de, 'h103df, 'h103e0, 'h103e1, 'h103e2, 'h103e3, 'h103e4, 'h103e5, 'h103e6, 'h103e7, 'h103e8, 'h103e9, 'h103ea, 'h103eb, 'h103ec, 'h103ed, 'h103ee, 'h103ef, 'h103f0, 'h103f1, 'h103f2, 'h103f3, 'h103f4, 'h103f5, 'h103f6, 'h103f7, 'h103f8, 'h103f9, 'h103fa, 'h103fb, 'h103fc, 'h103fd, 'h103fe, 'h103ff, 'h10400, 'h10401, 'h10402, 'h10403, 'h10404, 'h10405, 'h10406, 'h10407, 'h10408, 'h10409, 'h1040a, 'h1040b, 'h1040c, 'h1040d, 'h1040e, 'h1040f, 'h10410, 'h10411, 'h10412, 'h10413, 'h10414, 'h10415, 'h10416, 'h10417, 'h10418, 'h10419, 'h1041a, 'h1041b, 'h1041c, 'h1041d, 'h1041e, 'h1041f, 'h10420, 'h10421, 'h10422, 'h10423, 'h10424, 'h10425, 'h10426, 'h10427, 'h10428, 'h10429, 'h1042a, 'h1042b, 'h1042c, 'h1042d, 'h1042e, 'h1042f, 'h10430, 'h10431, 'h10432, 'h10433, 'h10434, 'h10435, 'h10436, 'h10437, 'h10438, 'h10439, 'h1043a, 'h1043b, 'h1043c, 'h1043d, 'h1043e, 'h1043f, 'h10442, 'h21f8c, 'h21f8a, 'h21f8b, 'h21f8d, 'h21f8f};
	
	int MM32_DATA [MM32_DATA_SIZE-1:0] = {DATA7, DATA0};
	
endpackage