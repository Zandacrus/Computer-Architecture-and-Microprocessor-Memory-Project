

package MATRIX_MULTIPLY_32_PKG_7;
	
	import MATRIX_MULTIPLY_32_PKG_6::DATA6;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h10849, 'h10ac9, 'h10cc9, 'h10859, 'h10869, 'h10aca, 'h10879, 'h10889, 'h10acb, 'h103bc, 'h10899, 'h108a9, 'h10acc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b9, 'h108c9, 'h10acd, 'h108d9, 'h106e9, 'h10ace, 'h10cd9, 'h106f9, 'h10709, 'h10acf, 'h10719, 'h10729, 'h10ad0, 'h10739, 'h103bc, 'h10749, 'h10ad1, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h10769, 'h10ad2, 'h10779, 'h10789, 'h10ad3, 'h10799, 'h10cd9, 'h107a9, 'h10ad4, 'h107b9, 'h107c9, 'h10ad5, 'h107d9, 'h107e9, 'h10ad6, 'h103bc, 'h107f9, 'h10809, 'h10ad7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10819, 'h10829, 'h10ad8, 'h10839, 'h10849, 'h10ad9, 'h10cd9, 'h10859, 'h10869, 'h10ada, 'h10879, 'h10889, 'h10adb, 'h10899, 'h103bc, 'h108a9, 'h10adc, 'h108b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c9, 'h10add, 'h108d9, 'h106ea, 'h108de, 'h10aea, 'h106fa, 'h1070a, 'h108df, 'h1071a, 'h1072a, 'h108e0, 'h1073a, 'h1074a, 'h108e1, 'h103bc, 'h1075a, 'h1076a, 'h108e2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077a, 'h1078a, 'h108e3, 'h1079a, 'h10aea, 'h107aa, 'h108e4, 'h107ba, 'h107ca, 'h108e5, 'h107da, 'h107ea, 'h108e6, 'h107fa, 'h103bc, 'h1080a, 'h108e7, 'h1081a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082a, 'h108e8, 'h1083a, 'h1084a, 'h108e9, 'h10aea, 'h1085a, 'h1086a, 'h108ea, 'h1087a, 'h1088a, 'h108eb, 'h1089a, 'h108aa, 'h108ec, 'h103bc, 'h108ba, 'h108ca, 'h108ed, 'h21f8e, 'h21f8f, 'h21f8d, 'h108da, 'h106ea, 'h108ee, 'h10afa, 'h106fa, 'h1070a, 'h108ef, 'h1071a, 'h1072a, 'h108f0, 'h1073a, 'h1074a, 'h108f1, 'h1075a, 'h103bc, 'h1076a, 'h108f2, 'h1077a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078a, 'h108f3, 'h1079a, 'h10afa, 'h107aa, 'h108f4, 'h107ba, 'h107ca, 'h108f5, 'h107da, 'h107ea, 'h108f6, 'h107fa, 'h1080a, 'h108f7, 'h103bc, 'h1081a, 'h1082a, 'h108f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083a, 'h1084a, 'h108f9, 'h10afa, 'h1085a, 'h1086a, 'h108fa, 'h1087a, 'h1088a, 'h108fb, 'h1089a, 'h108aa, 'h108fc, 'h108ba, 'h103bc, 'h108ca, 'h108fd, 'h108da, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ea, 'h108fe, 'h10b0a, 'h106fa, 'h1070a, 'h108ff, 'h1071a, 'h1072a, 'h10900, 'h1073a, 'h1074a, 'h10901, 'h1075a, 'h1076a, 'h10902, 'h103bc, 'h1077a, 'h1078a, 'h10903, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079a, 'h10b0a, 'h107aa, 'h10904, 'h107ba, 'h107ca, 'h10905, 'h107da, 'h107ea, 'h10906, 'h107fa, 'h1080a, 'h10907, 'h1081a, 'h103bc, 'h1082a, 'h10908, 'h1083a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084a, 'h10909, 'h10b0a, 'h1085a, 'h1086a, 'h1090a, 'h1087a, 'h1088a, 'h1090b, 'h1089a, 'h108aa, 'h1090c, 'h108ba, 'h108ca, 'h1090d, 'h103bc, 'h108da, 'h106ea, 'h1090e, 'h10b1a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fa, 'h1070a, 'h1090f, 'h1071a, 'h1072a, 'h10910, 'h1073a, 'h1074a, 'h10911, 'h1075a, 'h1076a, 'h10912, 'h1077a, 'h103bc, 'h1078a, 'h10913, 'h1079a, 'h10b1a, 'h21f8e, 'h21f8f, 'h21f8d, 'h107aa, 'h10914, 'h107ba, 'h107ca, 'h10915, 'h107da, 'h107ea, 'h10916, 'h107fa, 'h1080a, 'h10917, 'h1081a, 'h1082a, 'h10918, 'h103bc, 'h1083a, 'h1084a, 'h10919, 'h10b1a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085a, 'h1086a, 'h1091a, 'h1087a, 'h1088a, 'h1091b, 'h1089a, 'h108aa, 'h1091c, 'h108ba, 'h108ca, 'h1091d, 'h108da, 'h103bc, 'h106ea, 'h1091e, 'h10b2a, 'h106fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h1091f, 'h1071a, 'h1072a, 'h10920, 'h1073a, 'h1074a, 'h10921, 'h1075a, 'h1076a, 'h10922, 'h1077a, 'h1078a, 'h10923, 'h103bc, 'h1079a, 'h10b2a, 'h107aa, 'h10924, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ba, 'h107ca, 'h10925, 'h107da, 'h107ea, 'h10926, 'h107fa, 'h1080a, 'h10927, 'h1081a, 'h1082a, 'h10928, 'h1083a, 'h103bc, 'h1084a, 'h10929, 'h10b2a, 'h1085a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086a, 'h1092a, 'h1087a, 'h1088a, 'h1092b, 'h1089a, 'h108aa, 'h1092c, 'h108ba, 'h108ca, 'h1092d, 'h108da, 'h106ea, 'h1092e, 'h10b3a, 'h103bc, 'h106fa, 'h1070a, 'h1092f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071a, 'h1072a, 'h10930, 'h1073a, 'h1074a, 'h10931, 'h1075a, 'h1076a, 'h10932, 'h1077a, 'h1078a, 'h10933, 'h1079a, 'h10b3a, 'h103bc, 'h107aa, 'h10934, 'h107ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ca, 'h10935, 'h107da, 'h107ea, 'h10936, 'h107fa, 'h1080a, 'h10937, 'h1081a, 'h1082a, 'h10938, 'h1083a, 'h1084a, 'h10939, 'h10b3a, 'h103bc, 'h1085a, 'h1086a, 'h1093a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087a, 'h1088a, 'h1093b, 'h1089a, 'h108aa, 'h1093c, 'h108ba, 'h108ca, 'h1093d, 'h108da, 'h106ea, 'h1093e, 'h10b4a, 'h106fa, 'h103bc, 'h1070a, 'h1093f, 'h1071a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072a, 'h10940, 'h1073a, 'h1074a, 'h10941, 'h1075a, 'h1076a, 'h10942, 'h1077a, 'h1078a, 'h10943, 'h1079a, 'h10b4a, 'h107aa, 'h10944, 'h103bc, 'h107ba, 'h107ca, 'h10945, 'h21f8e, 'h21f8f, 'h21f8d, 'h107da, 'h107ea, 'h10946, 'h107fa, 'h1080a, 'h10947, 'h1081a, 'h1082a, 'h10948, 'h1083a, 'h1084a, 'h10949, 'h10b4a, 'h1085a, 'h103bc, 'h1086a, 'h1094a, 'h1087a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088a, 'h1094b, 'h1089a, 'h108aa, 'h1094c, 'h108ba, 'h108ca, 'h1094d, 'h108da, 'h106ea, 'h1094e, 'h10b5a, 'h106fa, 'h1070a, 'h1094f, 'h103bc, 'h1071a, 'h1072a, 'h10950, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h1074a, 'h10951, 'h1075a, 'h1076a, 'h10952, 'h1077a, 'h1078a, 'h10953, 'h1079a, 'h10b5a, 'h107aa, 'h10954, 'h107ba, 'h103bc, 'h107ca, 'h10955, 'h107da, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ea, 'h10956, 'h107fa, 'h1080a, 'h10957, 'h1081a, 'h1082a, 'h10958, 'h1083a, 'h1084a, 'h10959, 'h10b5a, 'h1085a, 'h1086a, 'h1095a, 'h103bc, 'h1087a, 'h1088a, 'h1095b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089a, 'h108aa, 'h1095c, 'h108ba, 'h108ca, 'h1095d, 'h108da, 'h106ea, 'h1095e, 'h10b6a, 'h106fa, 'h1070a, 'h1095f, 'h1071a, 'h103bc, 'h1072a, 'h10960, 'h1073a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074a, 'h10961, 'h1075a, 'h1076a, 'h10962, 'h1077a, 'h1078a, 'h10963, 'h1079a, 'h10b6a, 'h107aa, 'h10964, 'h107ba, 'h107ca, 'h10965, 'h103bc, 'h107da, 'h107ea, 'h10966, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fa, 'h1080a, 'h10967, 'h1081a, 'h1082a, 'h10968, 'h1083a, 'h1084a, 'h10969, 'h10b6a, 'h1085a, 'h1086a, 'h1096a, 'h1087a, 'h103bc, 'h1088a, 'h1096b, 'h1089a, 'h21f8e, 'h21f8f, 'h21f8d, 'h108aa, 'h1096c, 'h108ba, 'h108ca, 'h1096d, 'h108da, 'h106ea, 'h1096e, 'h10b7a, 'h106fa, 'h1070a, 'h1096f, 'h1071a, 'h1072a, 'h10970, 'h103bc, 'h1073a, 'h1074a, 'h10971, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075a, 'h1076a, 'h10972, 'h1077a, 'h1078a, 'h10973, 'h1079a, 'h10b7a, 'h107aa, 'h10974, 'h107ba, 'h107ca, 'h10975, 'h107da, 'h103bc, 'h107ea, 'h10976, 'h107fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080a, 'h10977, 'h1081a, 'h1082a, 'h10978, 'h1083a, 'h1084a, 'h10979, 'h10b7a, 'h1085a, 'h1086a, 'h1097a, 'h1087a, 'h1088a, 'h1097b, 'h103bc, 'h1089a, 'h108aa, 'h1097c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ba, 'h108ca, 'h1097d, 'h108da, 'h106ea, 'h1097e, 'h10b8a, 'h106fa, 'h1070a, 'h1097f, 'h1071a, 'h1072a, 'h10980, 'h1073a, 'h103bc, 'h1074a, 'h10981, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076a, 'h10982, 'h1077a, 'h1078a, 'h10983, 'h1079a, 'h10b8a, 'h107aa, 'h10984, 'h107ba, 'h107ca, 'h10985, 'h107da, 'h107ea, 'h10986, 'h103bc, 'h107fa, 'h1080a, 'h10987, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081a, 'h1082a, 'h10988, 'h1083a, 'h1084a, 'h10989, 'h10b8a, 'h1085a, 'h1086a, 'h1098a, 'h1087a, 'h1088a, 'h1098b, 'h1089a, 'h103bc, 'h108aa, 'h1098c, 'h108ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ca, 'h1098d, 'h108da, 'h106ea, 'h1098e, 'h10b9a, 'h106fa, 'h1070a, 'h1098f, 'h1071a, 'h1072a, 'h10990, 'h1073a, 'h1074a, 'h10991, 'h103bc, 'h1075a, 'h1076a, 'h10992, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077a, 'h1078a, 'h10993, 'h1079a, 'h10b9a, 'h107aa, 'h10994, 'h107ba, 'h107ca, 'h10995, 'h107da, 'h107ea, 'h10996, 'h107fa, 'h103bc, 'h1080a, 'h10997, 'h1081a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082a, 'h10998, 'h1083a, 'h1084a, 'h10999, 'h10b9a, 'h1085a, 'h1086a, 'h1099a, 'h1087a, 'h1088a, 'h1099b, 'h1089a, 'h108aa, 'h1099c, 'h103bc, 'h108ba, 'h108ca, 'h1099d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108da, 'h106ea, 'h1099e, 'h10baa, 'h106fa, 'h1070a, 'h1099f, 'h1071a, 'h1072a, 'h109a0, 'h1073a, 'h1074a, 'h109a1, 'h1075a, 'h103bc, 'h1076a, 'h109a2, 'h1077a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078a, 'h109a3, 'h1079a, 'h10baa, 'h107aa, 'h109a4, 'h107ba, 'h107ca, 'h109a5, 'h107da, 'h107ea, 'h109a6, 'h107fa, 'h1080a, 'h109a7, 'h103bc, 'h1081a, 'h1082a, 'h109a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083a, 'h1084a, 'h109a9, 'h10baa, 'h1085a, 'h1086a, 'h109aa, 'h1087a, 'h1088a, 'h109ab, 'h1089a, 'h108aa, 'h109ac, 'h108ba, 'h103bc, 'h108ca, 'h109ad, 'h108da, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ea, 'h109ae, 'h10bba, 'h106fa, 'h1070a, 'h109af, 'h1071a, 'h1072a, 'h109b0, 'h1073a, 'h1074a, 'h109b1, 'h1075a, 'h1076a, 'h109b2, 'h103bc, 'h1077a, 'h1078a, 'h109b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079a, 'h10bba, 'h107aa, 'h109b4, 'h107ba, 'h107ca, 'h109b5, 'h107da, 'h107ea, 'h109b6, 'h107fa, 'h1080a, 'h109b7, 'h1081a, 'h103bc, 'h1082a, 'h109b8, 'h1083a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084a, 'h109b9, 'h10bba, 'h1085a, 'h1086a, 'h109ba, 'h1087a, 'h1088a, 'h109bb, 'h1089a, 'h108aa, 'h109bc, 'h108ba, 'h108ca, 'h109bd, 'h103bc, 'h108da, 'h106ea, 'h109be, 'h10bca, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fa, 'h1070a, 'h109bf, 'h1071a, 'h1072a, 'h109c0, 'h1073a, 'h1074a, 'h109c1, 'h1075a, 'h1076a, 'h109c2, 'h1077a, 'h103bc, 'h1078a, 'h109c3, 'h1079a, 'h10bca, 'h21f8e, 'h21f8f, 'h21f8d, 'h107aa, 'h109c4, 'h107ba, 'h107ca, 'h109c5, 'h107da, 'h107ea, 'h109c6, 'h107fa, 'h1080a, 'h109c7, 'h1081a, 'h1082a, 'h109c8, 'h103bc, 'h1083a, 'h1084a, 'h109c9, 'h10bca, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085a, 'h1086a, 'h109ca, 'h1087a, 'h1088a, 'h109cb, 'h1089a, 'h108aa, 'h109cc, 'h108ba, 'h108ca, 'h109cd, 'h108da, 'h103bc, 'h106ea, 'h109ce, 'h10bda, 'h106fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h109cf, 'h1071a, 'h1072a, 'h109d0, 'h1073a, 'h1074a, 'h109d1, 'h1075a, 'h1076a, 'h109d2, 'h1077a, 'h1078a, 'h109d3, 'h103bc, 'h1079a, 'h10bda, 'h107aa, 'h109d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ba, 'h107ca, 'h109d5, 'h107da, 'h107ea, 'h109d6, 'h107fa, 'h1080a, 'h109d7, 'h1081a, 'h1082a, 'h109d8, 'h1083a, 'h103bc, 'h1084a, 'h109d9, 'h10bda, 'h1085a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086a, 'h109da, 'h1087a, 'h1088a, 'h109db, 'h1089a, 'h108aa, 'h109dc, 'h108ba, 'h108ca, 'h109dd, 'h108da, 'h106ea, 'h109de, 'h10bea, 'h103bc, 'h106fa, 'h1070a, 'h109df, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071a, 'h1072a, 'h109e0, 'h1073a, 'h1074a, 'h109e1, 'h1075a, 'h1076a, 'h109e2, 'h1077a, 'h1078a, 'h109e3, 'h1079a, 'h10bea, 'h103bc, 'h107aa, 'h109e4, 'h107ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ca, 'h109e5, 'h107da, 'h107ea, 'h109e6, 'h107fa, 'h1080a, 'h109e7, 'h1081a, 'h1082a, 'h109e8, 'h1083a, 'h1084a, 'h109e9, 'h10bea, 'h103bc, 'h1085a, 'h1086a, 'h109ea, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087a, 'h1088a, 'h109eb, 'h1089a, 'h108aa, 'h109ec, 'h108ba, 'h108ca, 'h109ed, 'h108da, 'h106ea, 'h109ee, 'h10bfa, 'h106fa, 'h103bc, 'h1070a, 'h109ef, 'h1071a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072a, 'h109f0, 'h1073a, 'h1074a, 'h109f1, 'h1075a, 'h1076a, 'h109f2, 'h1077a, 'h1078a, 'h109f3, 'h1079a, 'h10bfa, 'h107aa, 'h109f4, 'h103bc, 'h107ba, 'h107ca, 'h109f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107da, 'h107ea, 'h109f6, 'h107fa, 'h1080a, 'h109f7, 'h1081a, 'h1082a, 'h109f8, 'h1083a, 'h1084a, 'h109f9, 'h10bfa, 'h1085a, 'h103bc, 'h1086a, 'h109fa, 'h1087a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088a, 'h109fb, 'h1089a, 'h108aa, 'h109fc, 'h108ba, 'h108ca, 'h109fd, 'h108da, 'h106ea, 'h109fe, 'h10c0a, 'h106fa, 'h1070a, 'h109ff, 'h103bc, 'h1071a, 'h1072a, 'h10a00, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h1074a, 'h10a01, 'h1075a, 'h1076a, 'h10a02, 'h1077a, 'h1078a, 'h10a03, 'h1079a, 'h10c0a, 'h107aa, 'h10a04, 'h107ba, 'h103bc, 'h107ca, 'h10a05, 'h107da, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ea, 'h10a06, 'h107fa, 'h1080a, 'h10a07, 'h1081a, 'h1082a, 'h10a08, 'h1083a, 'h1084a, 'h10a09, 'h10c0a, 'h1085a, 'h1086a, 'h10a0a, 'h103bc, 'h1087a, 'h1088a, 'h10a0b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089a, 'h108aa, 'h10a0c, 'h108ba, 'h108ca, 'h10a0d, 'h108da, 'h106ea, 'h10a0e, 'h10c1a, 'h106fa, 'h1070a, 'h10a0f, 'h1071a, 'h103bc, 'h1072a, 'h10a10, 'h1073a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074a, 'h10a11, 'h1075a, 'h1076a, 'h10a12, 'h1077a, 'h1078a, 'h10a13, 'h1079a, 'h10c1a, 'h107aa, 'h10a14, 'h107ba, 'h107ca, 'h10a15, 'h103bc, 'h107da, 'h107ea, 'h10a16, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fa, 'h1080a, 'h10a17, 'h1081a, 'h1082a, 'h10a18, 'h1083a, 'h1084a, 'h10a19, 'h10c1a, 'h1085a, 'h1086a, 'h10a1a, 'h1087a, 'h103bc, 'h1088a, 'h10a1b, 'h1089a, 'h21f8e, 'h21f8f, 'h21f8d, 'h108aa, 'h10a1c, 'h108ba, 'h108ca, 'h10a1d, 'h108da, 'h106ea, 'h10a1e, 'h10c2a, 'h106fa, 'h1070a, 'h10a1f, 'h1071a, 'h1072a, 'h10a20, 'h103bc, 'h1073a, 'h1074a, 'h10a21, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075a, 'h1076a, 'h10a22, 'h1077a, 'h1078a, 'h10a23, 'h1079a, 'h10c2a, 'h107aa, 'h10a24, 'h107ba, 'h107ca, 'h10a25, 'h107da, 'h103bc, 'h107ea, 'h10a26, 'h107fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080a, 'h10a27, 'h1081a, 'h1082a, 'h10a28, 'h1083a, 'h1084a, 'h10a29, 'h10c2a, 'h1085a, 'h1086a, 'h10a2a, 'h1087a, 'h1088a, 'h10a2b, 'h103bc, 'h1089a, 'h108aa, 'h10a2c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ba, 'h108ca, 'h10a2d, 'h108da, 'h106ea, 'h10a2e, 'h10c3a, 'h106fa, 'h1070a, 'h10a2f, 'h1071a, 'h1072a, 'h10a30, 'h1073a, 'h103bc, 'h1074a, 'h10a31, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076a, 'h10a32, 'h1077a, 'h1078a, 'h10a33, 'h1079a, 'h10c3a, 'h107aa, 'h10a34, 'h107ba, 'h107ca, 'h10a35, 'h107da, 'h107ea, 'h10a36, 'h103bc, 'h107fa, 'h1080a, 'h10a37, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081a, 'h1082a, 'h10a38, 'h1083a, 'h1084a, 'h10a39, 'h10c3a, 'h1085a, 'h1086a, 'h10a3a, 'h1087a, 'h1088a, 'h10a3b, 'h1089a, 'h103bc, 'h108aa, 'h10a3c, 'h108ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ca, 'h10a3d, 'h108da, 'h106ea, 'h10a3e, 'h10c4a, 'h106fa, 'h1070a, 'h10a3f, 'h1071a, 'h1072a, 'h10a40, 'h1073a, 'h1074a, 'h10a41, 'h103bc, 'h1075a, 'h1076a, 'h10a42, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077a, 'h1078a, 'h10a43, 'h1079a, 'h10c4a, 'h107aa, 'h10a44, 'h107ba, 'h107ca, 'h10a45, 'h107da, 'h107ea, 'h10a46, 'h107fa, 'h103bc, 'h1080a, 'h10a47, 'h1081a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082a, 'h10a48, 'h1083a, 'h1084a, 'h10a49, 'h10c4a, 'h1085a, 'h1086a, 'h10a4a, 'h1087a, 'h1088a, 'h10a4b, 'h1089a, 'h108aa, 'h10a4c, 'h103bc, 'h108ba, 'h108ca, 'h10a4d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108da, 'h106ea, 'h10a4e, 'h10c5a, 'h106fa, 'h1070a, 'h10a4f, 'h1071a, 'h1072a, 'h10a50, 'h1073a, 'h1074a, 'h10a51, 'h1075a, 'h103bc, 'h1076a, 'h10a52, 'h1077a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078a, 'h10a53, 'h1079a, 'h10c5a, 'h107aa, 'h10a54, 'h107ba, 'h107ca, 'h10a55, 'h107da, 'h107ea, 'h10a56, 'h107fa, 'h1080a, 'h10a57, 'h103bc, 'h1081a, 'h1082a, 'h10a58, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083a, 'h1084a, 'h10a59, 'h10c5a, 'h1085a, 'h1086a, 'h10a5a, 'h1087a, 'h1088a, 'h10a5b, 'h1089a, 'h108aa, 'h10a5c, 'h108ba, 'h103bc, 'h108ca, 'h10a5d, 'h108da, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ea, 'h10a5e, 'h10c6a, 'h106fa, 'h1070a, 'h10a5f, 'h1071a, 'h1072a, 'h10a60, 'h1073a, 'h1074a, 'h10a61, 'h1075a, 'h1076a, 'h10a62, 'h103bc, 'h1077a, 'h1078a, 'h10a63, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079a, 'h10c6a, 'h107aa, 'h10a64, 'h107ba, 'h107ca, 'h10a65, 'h107da, 'h107ea, 'h10a66, 'h107fa, 'h1080a, 'h10a67, 'h1081a, 'h103bc, 'h1082a, 'h10a68, 'h1083a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084a, 'h10a69, 'h10c6a, 'h1085a, 'h1086a, 'h10a6a, 'h1087a, 'h1088a, 'h10a6b, 'h1089a, 'h108aa, 'h10a6c, 'h108ba, 'h108ca, 'h10a6d, 'h103bc, 'h108da, 'h106ea, 'h10a6e, 'h10c7a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fa, 'h1070a, 'h10a6f, 'h1071a, 'h1072a, 'h10a70, 'h1073a, 'h1074a, 'h10a71, 'h1075a, 'h1076a, 'h10a72, 'h1077a, 'h103bc, 'h1078a, 'h10a73, 'h1079a, 'h10c7a, 'h21f8e, 'h21f8f, 'h21f8d, 'h107aa, 'h10a74, 'h107ba, 'h107ca, 'h10a75, 'h107da, 'h107ea, 'h10a76, 'h107fa, 'h1080a, 'h10a77, 'h1081a, 'h1082a, 'h10a78, 'h103bc, 'h1083a, 'h1084a, 'h10a79, 'h10c7a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085a, 'h1086a, 'h10a7a, 'h1087a, 'h1088a, 'h10a7b, 'h1089a, 'h108aa, 'h10a7c, 'h108ba, 'h108ca, 'h10a7d, 'h108da, 'h103bc, 'h106ea, 'h10a7e, 'h10c8a, 'h106fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10a7f, 'h1071a, 'h1072a, 'h10a80, 'h1073a, 'h1074a, 'h10a81, 'h1075a, 'h1076a, 'h10a82, 'h1077a, 'h1078a, 'h10a83, 'h103bc, 'h1079a, 'h10c8a, 'h107aa, 'h10a84, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ba, 'h107ca, 'h10a85, 'h107da, 'h107ea, 'h10a86, 'h107fa, 'h1080a, 'h10a87, 'h1081a, 'h1082a, 'h10a88, 'h1083a, 'h103bc, 'h1084a, 'h10a89, 'h10c8a, 'h1085a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086a, 'h10a8a, 'h1087a, 'h1088a, 'h10a8b, 'h1089a, 'h108aa, 'h10a8c, 'h108ba, 'h108ca, 'h10a8d, 'h108da, 'h106ea, 'h10a8e, 'h10c9a, 'h103bc, 'h106fa, 'h1070a, 'h10a8f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071a, 'h1072a, 'h10a90, 'h1073a, 'h1074a, 'h10a91, 'h1075a, 'h1076a, 'h10a92, 'h1077a, 'h1078a, 'h10a93, 'h1079a, 'h10c9a, 'h103bc, 'h107aa, 'h10a94, 'h107ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ca, 'h10a95, 'h107da, 'h107ea, 'h10a96, 'h107fa, 'h1080a, 'h10a97, 'h1081a, 'h1082a, 'h10a98, 'h1083a, 'h1084a, 'h10a99, 'h10c9a, 'h103bc, 'h1085a, 'h1086a, 'h10a9a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087a, 'h1088a, 'h10a9b, 'h1089a, 'h108aa, 'h10a9c, 'h108ba, 'h108ca, 'h10a9d, 'h108da, 'h106ea, 'h10a9e, 'h10caa, 'h106fa, 'h103bc, 'h1070a, 'h10a9f, 'h1071a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072a, 'h10aa0, 'h1073a, 'h1074a, 'h10aa1, 'h1075a, 'h1076a, 'h10aa2, 'h1077a, 'h1078a, 'h10aa3, 'h1079a, 'h10caa, 'h107aa, 'h10aa4, 'h103bc, 'h107ba, 'h107ca, 'h10aa5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107da, 'h107ea, 'h10aa6, 'h107fa, 'h1080a, 'h10aa7, 'h1081a, 'h1082a, 'h10aa8, 'h1083a, 'h1084a, 'h10aa9, 'h10caa, 'h1085a, 'h103bc, 'h1086a, 'h10aaa, 'h1087a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088a, 'h10aab, 'h1089a, 'h108aa, 'h10aac, 'h108ba, 'h108ca, 'h10aad, 'h108da, 'h106ea, 'h10aae, 'h10cba, 'h106fa, 'h1070a, 'h10aaf, 'h103bc, 'h1071a, 'h1072a, 'h10ab0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h1074a, 'h10ab1, 'h1075a, 'h1076a, 'h10ab2, 'h1077a, 'h1078a, 'h10ab3, 'h1079a, 'h10cba, 'h107aa, 'h10ab4, 'h107ba, 'h103bc, 'h107ca, 'h10ab5, 'h107da, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ea, 'h10ab6, 'h107fa, 'h1080a, 'h10ab7, 'h1081a, 'h1082a, 'h10ab8, 'h1083a, 'h1084a, 'h10ab9, 'h10cba, 'h1085a, 'h1086a, 'h10aba, 'h103bc, 'h1087a, 'h1088a, 'h10abb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089a, 'h108aa, 'h10abc, 'h108ba, 'h108ca, 'h10abd, 'h108da, 'h106ea, 'h10abe, 'h10cca, 'h106fa, 'h1070a, 'h10abf, 'h1071a, 'h103bc, 'h1072a, 'h10ac0, 'h1073a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074a, 'h10ac1, 'h1075a, 'h1076a, 'h10ac2, 'h1077a, 'h1078a, 'h10ac3, 'h1079a, 'h10cca, 'h107aa, 'h10ac4, 'h107ba, 'h107ca, 'h10ac5, 'h103bc, 'h107da, 'h107ea, 'h10ac6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fa, 'h1080a, 'h10ac7, 'h1081a, 'h1082a, 'h10ac8, 'h1083a, 'h1084a, 'h10ac9, 'h10cca, 'h1085a, 'h1086a, 'h10aca, 'h1087a, 'h103bc, 'h1088a, 'h10acb, 'h1089a, 'h21f8e, 'h21f8f, 'h21f8d, 'h108aa, 'h10acc, 'h108ba, 'h108ca, 'h10acd, 'h108da, 'h106ea, 'h10ace, 'h10cda, 'h106fa, 'h1070a, 'h10acf, 'h1071a, 'h1072a, 'h10ad0, 'h103bc, 'h1073a, 'h1074a, 'h10ad1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075a, 'h1076a, 'h10ad2, 'h1077a, 'h1078a, 'h10ad3, 'h1079a, 'h10cda, 'h107aa, 'h10ad4, 'h107ba, 'h107ca, 'h10ad5, 'h107da, 'h103bc, 'h107ea, 'h10ad6, 'h107fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080a, 'h10ad7, 'h1081a, 'h1082a, 'h10ad8, 'h1083a, 'h1084a, 'h10ad9, 'h10cda, 'h1085a, 'h1086a, 'h10ada, 'h1087a, 'h1088a, 'h10adb, 'h103bc, 'h1089a, 'h108aa, 'h10adc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ba, 'h108ca, 'h10add, 'h108da, 'h106ea, 'h108de, 'h10aea, 'h106fa, 'h1070a, 'h108df, 'h1071a, 'h1072a, 'h108e0, 'h1073a, 'h103bc, 'h1074a, 'h108e1, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076a, 'h108e2, 'h1077a, 'h1078a, 'h108e3, 'h1079a, 'h10aea, 'h107aa, 'h108e4, 'h107ba, 'h107ca, 'h108e5, 'h107da, 'h107ea, 'h108e6, 'h103bc, 'h107fa, 'h1080a, 'h108e7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081a, 'h1082a, 'h108e8, 'h1083a, 'h1084a, 'h108e9, 'h10aea, 'h1085a, 'h1086a, 'h108ea, 'h1087a, 'h1088a, 'h108eb, 'h1089a, 'h103bc, 'h108aa, 'h108ec, 'h108ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ca, 'h108ed, 'h108da, 'h106ea, 'h108ee, 'h10afa, 'h106fa, 'h1070a, 'h108ef, 'h1071a, 'h1072a, 'h108f0, 'h1073a, 'h1074a, 'h108f1, 'h103bc, 'h1075a, 'h1076a, 'h108f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077a, 'h1078a, 'h108f3, 'h1079a, 'h10afa, 'h107aa, 'h108f4, 'h107ba, 'h107ca, 'h108f5, 'h107da, 'h107ea, 'h108f6, 'h107fa, 'h103bc, 'h1080a, 'h108f7, 'h1081a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082a, 'h108f8, 'h1083a, 'h1084a, 'h108f9, 'h10afa, 'h1085a, 'h1086a, 'h108fa, 'h1087a, 'h1088a, 'h108fb, 'h1089a, 'h108aa, 'h108fc, 'h103bc, 'h108ba, 'h108ca, 'h108fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108da, 'h106ea, 'h108fe, 'h10b0a, 'h106fa, 'h1070a, 'h108ff, 'h1071a, 'h1072a, 'h10900, 'h1073a, 'h1074a, 'h10901, 'h1075a, 'h103bc, 'h1076a, 'h10902, 'h1077a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078a, 'h10903, 'h1079a, 'h10b0a, 'h107aa, 'h10904, 'h107ba, 'h107ca, 'h10905, 'h107da, 'h107ea, 'h10906, 'h107fa, 'h1080a, 'h10907, 'h103bc, 'h1081a, 'h1082a, 'h10908, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083a, 'h1084a, 'h10909, 'h10b0a, 'h1085a, 'h1086a, 'h1090a, 'h1087a, 'h1088a, 'h1090b, 'h1089a, 'h108aa, 'h1090c, 'h108ba, 'h103bc, 'h108ca, 'h1090d, 'h108da, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ea, 'h1090e, 'h10b1a, 'h106fa, 'h1070a, 'h1090f, 'h1071a, 'h1072a, 'h10910, 'h1073a, 'h1074a, 'h10911, 'h1075a, 'h1076a, 'h10912, 'h103bc, 'h1077a, 'h1078a, 'h10913, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079a, 'h10b1a, 'h107aa, 'h10914, 'h107ba, 'h107ca, 'h10915, 'h107da, 'h107ea, 'h10916, 'h107fa, 'h1080a, 'h10917, 'h1081a, 'h103bc, 'h1082a, 'h10918, 'h1083a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084a, 'h10919, 'h10b1a, 'h1085a, 'h1086a, 'h1091a, 'h1087a, 'h1088a, 'h1091b, 'h1089a, 'h108aa, 'h1091c, 'h108ba, 'h108ca, 'h1091d, 'h103bc, 'h108da, 'h106ea, 'h1091e, 'h10b2a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fa, 'h1070a, 'h1091f, 'h1071a, 'h1072a, 'h10920, 'h1073a, 'h1074a, 'h10921, 'h1075a, 'h1076a, 'h10922, 'h1077a, 'h103bc, 'h1078a, 'h10923, 'h1079a, 'h10b2a, 'h21f8e, 'h21f8f, 'h21f8d, 'h107aa, 'h10924, 'h107ba, 'h107ca, 'h10925, 'h107da, 'h107ea, 'h10926, 'h107fa, 'h1080a, 'h10927, 'h1081a, 'h1082a, 'h10928, 'h103bc, 'h1083a, 'h1084a, 'h10929, 'h10b2a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085a, 'h1086a, 'h1092a, 'h1087a, 'h1088a, 'h1092b, 'h1089a, 'h108aa, 'h1092c, 'h108ba, 'h108ca, 'h1092d, 'h108da, 'h103bc, 'h106ea, 'h1092e, 'h10b3a, 'h106fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h1092f, 'h1071a, 'h1072a, 'h10930, 'h1073a, 'h1074a, 'h10931, 'h1075a, 'h1076a, 'h10932, 'h1077a, 'h1078a, 'h10933, 'h103bc, 'h1079a, 'h10b3a, 'h107aa, 'h10934, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ba, 'h107ca, 'h10935, 'h107da, 'h107ea, 'h10936, 'h107fa, 'h1080a, 'h10937, 'h1081a, 'h1082a, 'h10938, 'h1083a, 'h103bc, 'h1084a, 'h10939, 'h10b3a, 'h1085a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086a, 'h1093a, 'h1087a, 'h1088a, 'h1093b, 'h1089a, 'h108aa, 'h1093c, 'h108ba, 'h108ca, 'h1093d, 'h108da, 'h106ea, 'h1093e, 'h10b4a, 'h103bc, 'h106fa, 'h1070a, 'h1093f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071a, 'h1072a, 'h10940, 'h1073a, 'h1074a, 'h10941, 'h1075a, 'h1076a, 'h10942, 'h1077a, 'h1078a, 'h10943, 'h1079a, 'h10b4a, 'h103bc, 'h107aa, 'h10944, 'h107ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ca, 'h10945, 'h107da, 'h107ea, 'h10946, 'h107fa, 'h1080a, 'h10947, 'h1081a, 'h1082a, 'h10948, 'h1083a, 'h1084a, 'h10949, 'h10b4a, 'h103bc, 'h1085a, 'h1086a, 'h1094a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087a, 'h1088a, 'h1094b, 'h1089a, 'h108aa, 'h1094c, 'h108ba, 'h108ca, 'h1094d, 'h108da, 'h106ea, 'h1094e, 'h10b5a, 'h106fa, 'h103bc, 'h1070a, 'h1094f, 'h1071a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072a, 'h10950, 'h1073a, 'h1074a, 'h10951, 'h1075a, 'h1076a, 'h10952, 'h1077a, 'h1078a, 'h10953, 'h1079a, 'h10b5a, 'h107aa, 'h10954, 'h103bc, 'h107ba, 'h107ca, 'h10955, 'h21f8e, 'h21f8f, 'h21f8d, 'h107da, 'h107ea, 'h10956, 'h107fa, 'h1080a, 'h10957, 'h1081a, 'h1082a, 'h10958, 'h1083a, 'h1084a, 'h10959, 'h10b5a, 'h1085a, 'h103bc, 'h1086a, 'h1095a, 'h1087a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088a, 'h1095b, 'h1089a, 'h108aa, 'h1095c, 'h108ba, 'h108ca, 'h1095d, 'h108da, 'h106ea, 'h1095e, 'h10b6a, 'h106fa, 'h1070a, 'h1095f, 'h103bc, 'h1071a, 'h1072a, 'h10960, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h1074a, 'h10961, 'h1075a, 'h1076a, 'h10962, 'h1077a, 'h1078a, 'h10963, 'h1079a, 'h10b6a, 'h107aa, 'h10964, 'h107ba, 'h103bc, 'h107ca, 'h10965, 'h107da, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ea, 'h10966, 'h107fa, 'h1080a, 'h10967, 'h1081a, 'h1082a, 'h10968, 'h1083a, 'h1084a, 'h10969, 'h10b6a, 'h1085a, 'h1086a, 'h1096a, 'h103bc, 'h1087a, 'h1088a, 'h1096b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089a, 'h108aa, 'h1096c, 'h108ba, 'h108ca, 'h1096d, 'h108da, 'h106ea, 'h1096e, 'h10b7a, 'h106fa, 'h1070a, 'h1096f, 'h1071a, 'h103bc, 'h1072a, 'h10970, 'h1073a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074a, 'h10971, 'h1075a, 'h1076a, 'h10972, 'h1077a, 'h1078a, 'h10973, 'h1079a, 'h10b7a, 'h107aa, 'h10974, 'h107ba, 'h107ca, 'h10975, 'h103bc, 'h107da, 'h107ea, 'h10976, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fa, 'h1080a, 'h10977, 'h1081a, 'h1082a, 'h10978, 'h1083a, 'h1084a, 'h10979, 'h10b7a, 'h1085a, 'h1086a, 'h1097a, 'h1087a, 'h103bc, 'h1088a, 'h1097b, 'h1089a, 'h21f8e, 'h21f8f, 'h21f8d, 'h108aa, 'h1097c, 'h108ba, 'h108ca, 'h1097d, 'h108da, 'h106ea, 'h1097e, 'h10b8a, 'h106fa, 'h1070a, 'h1097f, 'h1071a, 'h1072a, 'h10980, 'h103bc, 'h1073a, 'h1074a, 'h10981, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075a, 'h1076a, 'h10982, 'h1077a, 'h1078a, 'h10983, 'h1079a, 'h10b8a, 'h107aa, 'h10984, 'h107ba, 'h107ca, 'h10985, 'h107da, 'h103bc, 'h107ea, 'h10986, 'h107fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080a, 'h10987, 'h1081a, 'h1082a, 'h10988, 'h1083a, 'h1084a, 'h10989, 'h10b8a, 'h1085a, 'h1086a, 'h1098a, 'h1087a, 'h1088a, 'h1098b, 'h103bc, 'h1089a, 'h108aa, 'h1098c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ba, 'h108ca, 'h1098d, 'h108da, 'h106ea, 'h1098e, 'h10b9a, 'h106fa, 'h1070a, 'h1098f, 'h1071a, 'h1072a, 'h10990, 'h1073a, 'h103bc, 'h1074a, 'h10991, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076a, 'h10992, 'h1077a, 'h1078a, 'h10993, 'h1079a, 'h10b9a, 'h107aa, 'h10994, 'h107ba, 'h107ca, 'h10995, 'h107da, 'h107ea, 'h10996, 'h103bc, 'h107fa, 'h1080a, 'h10997, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081a, 'h1082a, 'h10998, 'h1083a, 'h1084a, 'h10999, 'h10b9a, 'h1085a, 'h1086a, 'h1099a, 'h1087a, 'h1088a, 'h1099b, 'h1089a, 'h103bc, 'h108aa, 'h1099c, 'h108ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ca, 'h1099d, 'h108da, 'h106ea, 'h1099e, 'h10baa, 'h106fa, 'h1070a, 'h1099f, 'h1071a, 'h1072a, 'h109a0, 'h1073a, 'h1074a, 'h109a1, 'h103bc, 'h1075a, 'h1076a, 'h109a2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077a, 'h1078a, 'h109a3, 'h1079a, 'h10baa, 'h107aa, 'h109a4, 'h107ba, 'h107ca, 'h109a5, 'h107da, 'h107ea, 'h109a6, 'h107fa, 'h103bc, 'h1080a, 'h109a7, 'h1081a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082a, 'h109a8, 'h1083a, 'h1084a, 'h109a9, 'h10baa, 'h1085a, 'h1086a, 'h109aa, 'h1087a, 'h1088a, 'h109ab, 'h1089a, 'h108aa, 'h109ac, 'h103bc, 'h108ba, 'h108ca, 'h109ad, 'h21f8e, 'h21f8f, 'h21f8d, 'h108da, 'h106ea, 'h109ae, 'h10bba, 'h106fa, 'h1070a, 'h109af, 'h1071a, 'h1072a, 'h109b0, 'h1073a, 'h1074a, 'h109b1, 'h1075a, 'h103bc, 'h1076a, 'h109b2, 'h1077a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078a, 'h109b3, 'h1079a, 'h10bba, 'h107aa, 'h109b4, 'h107ba, 'h107ca, 'h109b5, 'h107da, 'h107ea, 'h109b6, 'h107fa, 'h1080a, 'h109b7, 'h103bc, 'h1081a, 'h1082a, 'h109b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083a, 'h1084a, 'h109b9, 'h10bba, 'h1085a, 'h1086a, 'h109ba, 'h1087a, 'h1088a, 'h109bb, 'h1089a, 'h108aa, 'h109bc, 'h108ba, 'h103bc, 'h108ca, 'h109bd, 'h108da, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ea, 'h109be, 'h10bca, 'h106fa, 'h1070a, 'h109bf, 'h1071a, 'h1072a, 'h109c0, 'h1073a, 'h1074a, 'h109c1, 'h1075a, 'h1076a, 'h109c2, 'h103bc, 'h1077a, 'h1078a, 'h109c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079a, 'h10bca, 'h107aa, 'h109c4, 'h107ba, 'h107ca, 'h109c5, 'h107da, 'h107ea, 'h109c6, 'h107fa, 'h1080a, 'h109c7, 'h1081a, 'h103bc, 'h1082a, 'h109c8, 'h1083a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084a, 'h109c9, 'h10bca, 'h1085a, 'h1086a, 'h109ca, 'h1087a, 'h1088a, 'h109cb, 'h1089a, 'h108aa, 'h109cc, 'h108ba, 'h108ca, 'h109cd, 'h103bc, 'h108da, 'h106ea, 'h109ce, 'h10bda, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fa, 'h1070a, 'h109cf, 'h1071a, 'h1072a, 'h109d0, 'h1073a, 'h1074a, 'h109d1, 'h1075a, 'h1076a, 'h109d2, 'h1077a, 'h103bc, 'h1078a, 'h109d3, 'h1079a, 'h10bda, 'h21f8e, 'h21f8f, 'h21f8d, 'h107aa, 'h109d4, 'h107ba, 'h107ca, 'h109d5, 'h107da, 'h107ea, 'h109d6, 'h107fa, 'h1080a, 'h109d7, 'h1081a, 'h1082a, 'h109d8, 'h103bc, 'h1083a, 'h1084a, 'h109d9, 'h10bda, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085a, 'h1086a, 'h109da, 'h1087a, 'h1088a, 'h109db, 'h1089a, 'h108aa, 'h109dc, 'h108ba, 'h108ca, 'h109dd, 'h108da, 'h103bc, 'h106ea, 'h109de, 'h10bea, 'h106fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h109df, 'h1071a, 'h1072a, 'h109e0, 'h1073a, 'h1074a, 'h109e1, 'h1075a, 'h1076a, 'h109e2, 'h1077a, 'h1078a, 'h109e3, 'h103bc, 'h1079a, 'h10bea, 'h107aa, 'h109e4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ba, 'h107ca, 'h109e5, 'h107da, 'h107ea, 'h109e6, 'h107fa, 'h1080a, 'h109e7, 'h1081a, 'h1082a, 'h109e8, 'h1083a, 'h103bc, 'h1084a, 'h109e9, 'h10bea, 'h1085a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086a, 'h109ea, 'h1087a, 'h1088a, 'h109eb, 'h1089a, 'h108aa, 'h109ec, 'h108ba, 'h108ca, 'h109ed, 'h108da, 'h106ea, 'h109ee, 'h10bfa, 'h103bc, 'h106fa, 'h1070a, 'h109ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071a, 'h1072a, 'h109f0, 'h1073a, 'h1074a, 'h109f1, 'h1075a, 'h1076a, 'h109f2, 'h1077a, 'h1078a, 'h109f3, 'h1079a, 'h10bfa, 'h103bc, 'h107aa, 'h109f4, 'h107ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ca, 'h109f5, 'h107da, 'h107ea, 'h109f6, 'h107fa, 'h1080a, 'h109f7, 'h1081a, 'h1082a, 'h109f8, 'h1083a, 'h1084a, 'h109f9, 'h10bfa, 'h103bc, 'h1085a, 'h1086a, 'h109fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087a, 'h1088a, 'h109fb, 'h1089a, 'h108aa, 'h109fc, 'h108ba, 'h108ca, 'h109fd, 'h108da, 'h106ea, 'h109fe, 'h10c0a, 'h106fa, 'h103bc, 'h1070a, 'h109ff, 'h1071a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072a, 'h10a00, 'h1073a, 'h1074a, 'h10a01, 'h1075a, 'h1076a, 'h10a02, 'h1077a, 'h1078a, 'h10a03, 'h1079a, 'h10c0a, 'h107aa, 'h10a04, 'h103bc, 'h107ba, 'h107ca, 'h10a05, 'h21f8e, 'h21f8f, 'h21f8d, 'h107da, 'h107ea, 'h10a06, 'h107fa, 'h1080a, 'h10a07, 'h1081a, 'h1082a, 'h10a08, 'h1083a, 'h1084a, 'h10a09, 'h10c0a, 'h1085a, 'h103bc, 'h1086a, 'h10a0a, 'h1087a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088a, 'h10a0b, 'h1089a, 'h108aa, 'h10a0c, 'h108ba, 'h108ca, 'h10a0d, 'h108da, 'h106ea, 'h10a0e, 'h10c1a, 'h106fa, 'h1070a, 'h10a0f, 'h103bc, 'h1071a, 'h1072a, 'h10a10, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h1074a, 'h10a11, 'h1075a, 'h1076a, 'h10a12, 'h1077a, 'h1078a, 'h10a13, 'h1079a, 'h10c1a, 'h107aa, 'h10a14, 'h107ba, 'h103bc, 'h107ca, 'h10a15, 'h107da, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ea, 'h10a16, 'h107fa, 'h1080a, 'h10a17, 'h1081a, 'h1082a, 'h10a18, 'h1083a, 'h1084a, 'h10a19, 'h10c1a, 'h1085a, 'h1086a, 'h10a1a, 'h103bc, 'h1087a, 'h1088a, 'h10a1b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089a, 'h108aa, 'h10a1c, 'h108ba, 'h108ca, 'h10a1d, 'h108da, 'h106ea, 'h10a1e, 'h10c2a, 'h106fa, 'h1070a, 'h10a1f, 'h1071a, 'h103bc, 'h1072a, 'h10a20, 'h1073a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074a, 'h10a21, 'h1075a, 'h1076a, 'h10a22, 'h1077a, 'h1078a, 'h10a23, 'h1079a, 'h10c2a, 'h107aa, 'h10a24, 'h107ba, 'h107ca, 'h10a25, 'h103bc, 'h107da, 'h107ea, 'h10a26, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fa, 'h1080a, 'h10a27, 'h1081a, 'h1082a, 'h10a28, 'h1083a, 'h1084a, 'h10a29, 'h10c2a, 'h1085a, 'h1086a, 'h10a2a, 'h1087a, 'h103bc, 'h1088a, 'h10a2b, 'h1089a, 'h21f8e, 'h21f8f, 'h21f8d, 'h108aa, 'h10a2c, 'h108ba, 'h108ca, 'h10a2d, 'h108da, 'h106ea, 'h10a2e, 'h10c3a, 'h106fa, 'h1070a, 'h10a2f, 'h1071a, 'h1072a, 'h10a30, 'h103bc, 'h1073a, 'h1074a, 'h10a31, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075a, 'h1076a, 'h10a32, 'h1077a, 'h1078a, 'h10a33, 'h1079a, 'h10c3a, 'h107aa, 'h10a34, 'h107ba, 'h107ca, 'h10a35, 'h107da, 'h103bc, 'h107ea, 'h10a36, 'h107fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080a, 'h10a37, 'h1081a, 'h1082a, 'h10a38, 'h1083a, 'h1084a, 'h10a39, 'h10c3a, 'h1085a, 'h1086a, 'h10a3a, 'h1087a, 'h1088a, 'h10a3b, 'h103bc, 'h1089a, 'h108aa, 'h10a3c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ba, 'h108ca, 'h10a3d, 'h108da, 'h106ea, 'h10a3e, 'h10c4a, 'h106fa, 'h1070a, 'h10a3f, 'h1071a, 'h1072a, 'h10a40, 'h1073a, 'h103bc, 'h1074a, 'h10a41, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076a, 'h10a42, 'h1077a, 'h1078a, 'h10a43, 'h1079a, 'h10c4a, 'h107aa, 'h10a44, 'h107ba, 'h107ca, 'h10a45, 'h107da, 'h107ea, 'h10a46, 'h103bc, 'h107fa, 'h1080a, 'h10a47, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081a, 'h1082a, 'h10a48, 'h1083a, 'h1084a, 'h10a49, 'h10c4a, 'h1085a, 'h1086a, 'h10a4a, 'h1087a, 'h1088a, 'h10a4b, 'h1089a, 'h103bc, 'h108aa, 'h10a4c, 'h108ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ca, 'h10a4d, 'h108da, 'h106ea, 'h10a4e, 'h10c5a, 'h106fa, 'h1070a, 'h10a4f, 'h1071a, 'h1072a, 'h10a50, 'h1073a, 'h1074a, 'h10a51, 'h103bc, 'h1075a, 'h1076a, 'h10a52, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077a, 'h1078a, 'h10a53, 'h1079a, 'h10c5a, 'h107aa, 'h10a54, 'h107ba, 'h107ca, 'h10a55, 'h107da, 'h107ea, 'h10a56, 'h107fa, 'h103bc, 'h1080a, 'h10a57, 'h1081a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082a, 'h10a58, 'h1083a, 'h1084a, 'h10a59, 'h10c5a, 'h1085a, 'h1086a, 'h10a5a, 'h1087a, 'h1088a, 'h10a5b, 'h1089a, 'h108aa, 'h10a5c, 'h103bc, 'h108ba, 'h108ca, 'h10a5d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108da, 'h106ea, 'h10a5e, 'h10c6a, 'h106fa, 'h1070a, 'h10a5f, 'h1071a, 'h1072a, 'h10a60, 'h1073a, 'h1074a, 'h10a61, 'h1075a, 'h103bc, 'h1076a, 'h10a62, 'h1077a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078a, 'h10a63, 'h1079a, 'h10c6a, 'h107aa, 'h10a64, 'h107ba, 'h107ca, 'h10a65, 'h107da, 'h107ea, 'h10a66, 'h107fa, 'h1080a, 'h10a67, 'h103bc, 'h1081a, 'h1082a, 'h10a68, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083a, 'h1084a, 'h10a69, 'h10c6a, 'h1085a, 'h1086a, 'h10a6a, 'h1087a, 'h1088a, 'h10a6b, 'h1089a, 'h108aa, 'h10a6c, 'h108ba, 'h103bc, 'h108ca, 'h10a6d, 'h108da, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ea, 'h10a6e, 'h10c7a, 'h106fa, 'h1070a, 'h10a6f, 'h1071a, 'h1072a, 'h10a70, 'h1073a, 'h1074a, 'h10a71, 'h1075a, 'h1076a, 'h10a72, 'h103bc, 'h1077a, 'h1078a, 'h10a73, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079a, 'h10c7a, 'h107aa, 'h10a74, 'h107ba, 'h107ca, 'h10a75, 'h107da, 'h107ea, 'h10a76, 'h107fa, 'h1080a, 'h10a77, 'h1081a, 'h103bc, 'h1082a, 'h10a78, 'h1083a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084a, 'h10a79, 'h10c7a, 'h1085a, 'h1086a, 'h10a7a, 'h1087a, 'h1088a, 'h10a7b, 'h1089a, 'h108aa, 'h10a7c, 'h108ba, 'h108ca, 'h10a7d, 'h103bc, 'h108da, 'h106ea, 'h10a7e, 'h10c8a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fa, 'h1070a, 'h10a7f, 'h1071a, 'h1072a, 'h10a80, 'h1073a, 'h1074a, 'h10a81, 'h1075a, 'h1076a, 'h10a82, 'h1077a, 'h103bc, 'h1078a, 'h10a83, 'h1079a, 'h10c8a, 'h21f8e, 'h21f8f, 'h21f8d, 'h107aa, 'h10a84, 'h107ba, 'h107ca, 'h10a85, 'h107da, 'h107ea, 'h10a86, 'h107fa, 'h1080a, 'h10a87, 'h1081a, 'h1082a, 'h10a88, 'h103bc, 'h1083a, 'h1084a, 'h10a89, 'h10c8a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085a, 'h1086a, 'h10a8a, 'h1087a, 'h1088a, 'h10a8b, 'h1089a, 'h108aa, 'h10a8c, 'h108ba, 'h108ca, 'h10a8d, 'h108da, 'h103bc, 'h106ea, 'h10a8e, 'h10c9a, 'h106fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10a8f, 'h1071a, 'h1072a, 'h10a90, 'h1073a, 'h1074a, 'h10a91, 'h1075a, 'h1076a, 'h10a92, 'h1077a, 'h1078a, 'h10a93, 'h103bc, 'h1079a, 'h10c9a, 'h107aa, 'h10a94, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ba, 'h107ca, 'h10a95, 'h107da, 'h107ea, 'h10a96, 'h107fa, 'h1080a, 'h10a97, 'h1081a, 'h1082a, 'h10a98, 'h1083a, 'h103bc, 'h1084a, 'h10a99, 'h10c9a, 'h1085a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086a, 'h10a9a, 'h1087a, 'h1088a, 'h10a9b, 'h1089a, 'h108aa, 'h10a9c, 'h108ba, 'h108ca, 'h10a9d, 'h108da, 'h106ea, 'h10a9e, 'h10caa, 'h103bc, 'h106fa, 'h1070a, 'h10a9f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071a, 'h1072a, 'h10aa0, 'h1073a, 'h1074a, 'h10aa1, 'h1075a, 'h1076a, 'h10aa2, 'h1077a, 'h1078a, 'h10aa3, 'h1079a, 'h10caa, 'h103bc, 'h107aa, 'h10aa4, 'h107ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ca, 'h10aa5, 'h107da, 'h107ea, 'h10aa6, 'h107fa, 'h1080a, 'h10aa7, 'h1081a, 'h1082a, 'h10aa8, 'h1083a, 'h1084a, 'h10aa9, 'h10caa, 'h103bc, 'h1085a, 'h1086a, 'h10aaa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087a, 'h1088a, 'h10aab, 'h1089a, 'h108aa, 'h10aac, 'h108ba, 'h108ca, 'h10aad, 'h108da, 'h106ea, 'h10aae, 'h10cba, 'h106fa, 'h103bc, 'h1070a, 'h10aaf, 'h1071a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072a, 'h10ab0, 'h1073a, 'h1074a, 'h10ab1, 'h1075a, 'h1076a, 'h10ab2, 'h1077a, 'h1078a, 'h10ab3, 'h1079a, 'h10cba, 'h107aa, 'h10ab4, 'h103bc, 'h107ba, 'h107ca, 'h10ab5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107da, 'h107ea, 'h10ab6, 'h107fa, 'h1080a, 'h10ab7, 'h1081a, 'h1082a, 'h10ab8, 'h1083a, 'h1084a, 'h10ab9, 'h10cba, 'h1085a, 'h103bc, 'h1086a, 'h10aba, 'h1087a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088a, 'h10abb, 'h1089a, 'h108aa, 'h10abc, 'h108ba, 'h108ca, 'h10abd, 'h108da, 'h106ea, 'h10abe, 'h10cca, 'h106fa, 'h1070a, 'h10abf, 'h103bc, 'h1071a, 'h1072a, 'h10ac0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h1074a, 'h10ac1, 'h1075a, 'h1076a, 'h10ac2, 'h1077a, 'h1078a, 'h10ac3, 'h1079a, 'h10cca, 'h107aa, 'h10ac4, 'h107ba, 'h103bc, 'h107ca, 'h10ac5, 'h107da, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ea, 'h10ac6, 'h107fa, 'h1080a, 'h10ac7, 'h1081a, 'h1082a, 'h10ac8, 'h1083a, 'h1084a, 'h10ac9, 'h10cca, 'h1085a, 'h1086a, 'h10aca, 'h103bc, 'h1087a, 'h1088a, 'h10acb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089a, 'h108aa, 'h10acc, 'h108ba, 'h108ca, 'h10acd, 'h108da, 'h106ea, 'h10ace, 'h10cda, 'h106fa, 'h1070a, 'h10acf, 'h1071a, 'h103bc, 'h1072a, 'h10ad0, 'h1073a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074a, 'h10ad1, 'h1075a, 'h1076a, 'h10ad2, 'h1077a, 'h1078a, 'h10ad3, 'h1079a, 'h10cda, 'h107aa, 'h10ad4, 'h107ba, 'h107ca, 'h10ad5, 'h103bc, 'h107da, 'h107ea, 'h10ad6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fa, 'h1080a, 'h10ad7, 'h1081a, 'h1082a, 'h10ad8, 'h1083a, 'h1084a, 'h10ad9, 'h10cda, 'h1085a, 'h1086a, 'h10ada, 'h1087a, 'h103bc, 'h1088a, 'h10adb, 'h1089a, 'h21f8e, 'h21f8f, 'h21f8d, 'h108aa, 'h10adc, 'h108ba, 'h108ca, 'h10add, 'h108da, 'h106eb, 'h108de, 'h10aeb, 'h106fb, 'h1070b, 'h108df, 'h1071b, 'h1072b, 'h108e0, 'h103bc, 'h1073b, 'h1074b, 'h108e1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075b, 'h1076b, 'h108e2, 'h1077b, 'h1078b, 'h108e3, 'h1079b, 'h10aeb, 'h107ab, 'h108e4, 'h107bb, 'h107cb, 'h108e5, 'h107db, 'h103bc, 'h107eb, 'h108e6, 'h107fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080b, 'h108e7, 'h1081b, 'h1082b, 'h108e8, 'h1083b, 'h1084b, 'h108e9, 'h10aeb, 'h1085b, 'h1086b, 'h108ea, 'h1087b, 'h1088b, 'h108eb, 'h103bc, 'h1089b, 'h108ab, 'h108ec, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bb, 'h108cb, 'h108ed, 'h108db, 'h106eb, 'h108ee, 'h10afb, 'h106fb, 'h1070b, 'h108ef, 'h1071b, 'h1072b, 'h108f0, 'h1073b, 'h103bc, 'h1074b, 'h108f1, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076b, 'h108f2, 'h1077b, 'h1078b, 'h108f3, 'h1079b, 'h10afb, 'h107ab, 'h108f4, 'h107bb, 'h107cb, 'h108f5, 'h107db, 'h107eb, 'h108f6, 'h103bc, 'h107fb, 'h1080b, 'h108f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081b, 'h1082b, 'h108f8, 'h1083b, 'h1084b, 'h108f9, 'h10afb, 'h1085b, 'h1086b, 'h108fa, 'h1087b, 'h1088b, 'h108fb, 'h1089b, 'h103bc, 'h108ab, 'h108fc, 'h108bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cb, 'h108fd, 'h108db, 'h106eb, 'h108fe, 'h10b0b, 'h106fb, 'h1070b, 'h108ff, 'h1071b, 'h1072b, 'h10900, 'h1073b, 'h1074b, 'h10901, 'h103bc, 'h1075b, 'h1076b, 'h10902, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077b, 'h1078b, 'h10903, 'h1079b, 'h10b0b, 'h107ab, 'h10904, 'h107bb, 'h107cb, 'h10905, 'h107db, 'h107eb, 'h10906, 'h107fb, 'h103bc, 'h1080b, 'h10907, 'h1081b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082b, 'h10908, 'h1083b, 'h1084b, 'h10909, 'h10b0b, 'h1085b, 'h1086b, 'h1090a, 'h1087b, 'h1088b, 'h1090b, 'h1089b, 'h108ab, 'h1090c, 'h103bc, 'h108bb, 'h108cb, 'h1090d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108db, 'h106eb, 'h1090e, 'h10b1b, 'h106fb, 'h1070b, 'h1090f, 'h1071b, 'h1072b, 'h10910, 'h1073b, 'h1074b, 'h10911, 'h1075b, 'h103bc, 'h1076b, 'h10912, 'h1077b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078b, 'h10913, 'h1079b, 'h10b1b, 'h107ab, 'h10914, 'h107bb, 'h107cb, 'h10915, 'h107db, 'h107eb, 'h10916, 'h107fb, 'h1080b, 'h10917, 'h103bc, 'h1081b, 'h1082b, 'h10918, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083b, 'h1084b, 'h10919, 'h10b1b, 'h1085b, 'h1086b, 'h1091a, 'h1087b, 'h1088b, 'h1091b, 'h1089b, 'h108ab, 'h1091c, 'h108bb, 'h103bc, 'h108cb, 'h1091d, 'h108db, 'h21f8e, 'h21f8f, 'h21f8d, 'h106eb, 'h1091e, 'h10b2b, 'h106fb, 'h1070b, 'h1091f, 'h1071b, 'h1072b, 'h10920, 'h1073b, 'h1074b, 'h10921, 'h1075b, 'h1076b, 'h10922, 'h103bc, 'h1077b, 'h1078b, 'h10923, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079b, 'h10b2b, 'h107ab, 'h10924, 'h107bb, 'h107cb, 'h10925, 'h107db, 'h107eb, 'h10926, 'h107fb, 'h1080b, 'h10927, 'h1081b, 'h103bc, 'h1082b, 'h10928, 'h1083b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084b, 'h10929, 'h10b2b, 'h1085b, 'h1086b, 'h1092a, 'h1087b, 'h1088b, 'h1092b, 'h1089b, 'h108ab, 'h1092c, 'h108bb, 'h108cb, 'h1092d, 'h103bc, 'h108db, 'h106eb, 'h1092e, 'h10b3b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fb, 'h1070b, 'h1092f, 'h1071b, 'h1072b, 'h10930, 'h1073b, 'h1074b, 'h10931, 'h1075b, 'h1076b, 'h10932, 'h1077b, 'h103bc, 'h1078b, 'h10933, 'h1079b, 'h10b3b, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ab, 'h10934, 'h107bb, 'h107cb, 'h10935, 'h107db, 'h107eb, 'h10936, 'h107fb, 'h1080b, 'h10937, 'h1081b, 'h1082b, 'h10938, 'h103bc, 'h1083b, 'h1084b, 'h10939, 'h10b3b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085b, 'h1086b, 'h1093a, 'h1087b, 'h1088b, 'h1093b, 'h1089b, 'h108ab, 'h1093c, 'h108bb, 'h108cb, 'h1093d, 'h108db, 'h103bc, 'h106eb, 'h1093e, 'h10b4b, 'h106fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h1093f, 'h1071b, 'h1072b, 'h10940, 'h1073b, 'h1074b, 'h10941, 'h1075b, 'h1076b, 'h10942, 'h1077b, 'h1078b, 'h10943, 'h103bc, 'h1079b, 'h10b4b, 'h107ab, 'h10944, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bb, 'h107cb, 'h10945, 'h107db, 'h107eb, 'h10946, 'h107fb, 'h1080b, 'h10947, 'h1081b, 'h1082b, 'h10948, 'h1083b, 'h103bc, 'h1084b, 'h10949, 'h10b4b, 'h1085b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086b, 'h1094a, 'h1087b, 'h1088b, 'h1094b, 'h1089b, 'h108ab, 'h1094c, 'h108bb, 'h108cb, 'h1094d, 'h108db, 'h106eb, 'h1094e, 'h10b5b, 'h103bc, 'h106fb, 'h1070b, 'h1094f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071b, 'h1072b, 'h10950, 'h1073b, 'h1074b, 'h10951, 'h1075b, 'h1076b, 'h10952, 'h1077b, 'h1078b, 'h10953, 'h1079b, 'h10b5b, 'h103bc, 'h107ab, 'h10954, 'h107bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cb, 'h10955, 'h107db, 'h107eb, 'h10956, 'h107fb, 'h1080b, 'h10957, 'h1081b, 'h1082b, 'h10958, 'h1083b, 'h1084b, 'h10959, 'h10b5b, 'h103bc, 'h1085b, 'h1086b, 'h1095a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087b, 'h1088b, 'h1095b, 'h1089b, 'h108ab, 'h1095c, 'h108bb, 'h108cb, 'h1095d, 'h108db, 'h106eb, 'h1095e, 'h10b6b, 'h106fb, 'h103bc, 'h1070b, 'h1095f, 'h1071b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072b, 'h10960, 'h1073b, 'h1074b, 'h10961, 'h1075b, 'h1076b, 'h10962, 'h1077b, 'h1078b, 'h10963, 'h1079b, 'h10b6b, 'h107ab, 'h10964, 'h103bc, 'h107bb, 'h107cb, 'h10965, 'h21f8e, 'h21f8f, 'h21f8d, 'h107db, 'h107eb, 'h10966, 'h107fb, 'h1080b, 'h10967, 'h1081b, 'h1082b, 'h10968, 'h1083b, 'h1084b, 'h10969, 'h10b6b, 'h1085b, 'h103bc, 'h1086b, 'h1096a, 'h1087b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088b, 'h1096b, 'h1089b, 'h108ab, 'h1096c, 'h108bb, 'h108cb, 'h1096d, 'h108db, 'h106eb, 'h1096e, 'h10b7b, 'h106fb, 'h1070b, 'h1096f, 'h103bc, 'h1071b, 'h1072b, 'h10970, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h1074b, 'h10971, 'h1075b, 'h1076b, 'h10972, 'h1077b, 'h1078b, 'h10973, 'h1079b, 'h10b7b, 'h107ab, 'h10974, 'h107bb, 'h103bc, 'h107cb, 'h10975, 'h107db, 'h21f8e, 'h21f8f, 'h21f8d, 'h107eb, 'h10976, 'h107fb, 'h1080b, 'h10977, 'h1081b, 'h1082b, 'h10978, 'h1083b, 'h1084b, 'h10979, 'h10b7b, 'h1085b, 'h1086b, 'h1097a, 'h103bc, 'h1087b, 'h1088b, 'h1097b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089b, 'h108ab, 'h1097c, 'h108bb, 'h108cb, 'h1097d, 'h108db, 'h106eb, 'h1097e, 'h10b8b, 'h106fb, 'h1070b, 'h1097f, 'h1071b, 'h103bc, 'h1072b, 'h10980, 'h1073b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074b, 'h10981, 'h1075b, 'h1076b, 'h10982, 'h1077b, 'h1078b, 'h10983, 'h1079b, 'h10b8b, 'h107ab, 'h10984, 'h107bb, 'h107cb, 'h10985, 'h103bc, 'h107db, 'h107eb, 'h10986, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fb, 'h1080b, 'h10987, 'h1081b, 'h1082b, 'h10988, 'h1083b, 'h1084b, 'h10989, 'h10b8b, 'h1085b, 'h1086b, 'h1098a, 'h1087b, 'h103bc, 'h1088b, 'h1098b, 'h1089b, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ab, 'h1098c, 'h108bb, 'h108cb, 'h1098d, 'h108db, 'h106eb, 'h1098e, 'h10b9b, 'h106fb, 'h1070b, 'h1098f, 'h1071b, 'h1072b, 'h10990, 'h103bc, 'h1073b, 'h1074b, 'h10991, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075b, 'h1076b, 'h10992, 'h1077b, 'h1078b, 'h10993, 'h1079b, 'h10b9b, 'h107ab, 'h10994, 'h107bb, 'h107cb, 'h10995, 'h107db, 'h103bc, 'h107eb, 'h10996, 'h107fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080b, 'h10997, 'h1081b, 'h1082b, 'h10998, 'h1083b, 'h1084b, 'h10999, 'h10b9b, 'h1085b, 'h1086b, 'h1099a, 'h1087b, 'h1088b, 'h1099b, 'h103bc, 'h1089b, 'h108ab, 'h1099c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bb, 'h108cb, 'h1099d, 'h108db, 'h106eb, 'h1099e, 'h10bab, 'h106fb, 'h1070b, 'h1099f, 'h1071b, 'h1072b, 'h109a0, 'h1073b, 'h103bc, 'h1074b, 'h109a1, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076b, 'h109a2, 'h1077b, 'h1078b, 'h109a3, 'h1079b, 'h10bab, 'h107ab, 'h109a4, 'h107bb, 'h107cb, 'h109a5, 'h107db, 'h107eb, 'h109a6, 'h103bc, 'h107fb, 'h1080b, 'h109a7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081b, 'h1082b, 'h109a8, 'h1083b, 'h1084b, 'h109a9, 'h10bab, 'h1085b, 'h1086b, 'h109aa, 'h1087b, 'h1088b, 'h109ab, 'h1089b, 'h103bc, 'h108ab, 'h109ac, 'h108bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cb, 'h109ad, 'h108db, 'h106eb, 'h109ae, 'h10bbb, 'h106fb, 'h1070b, 'h109af, 'h1071b, 'h1072b, 'h109b0, 'h1073b, 'h1074b, 'h109b1, 'h103bc, 'h1075b, 'h1076b, 'h109b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077b, 'h1078b, 'h109b3, 'h1079b, 'h10bbb, 'h107ab, 'h109b4, 'h107bb, 'h107cb, 'h109b5, 'h107db, 'h107eb, 'h109b6, 'h107fb, 'h103bc, 'h1080b, 'h109b7, 'h1081b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082b, 'h109b8, 'h1083b, 'h1084b, 'h109b9, 'h10bbb, 'h1085b, 'h1086b, 'h109ba, 'h1087b, 'h1088b, 'h109bb, 'h1089b, 'h108ab, 'h109bc, 'h103bc, 'h108bb, 'h108cb, 'h109bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108db, 'h106eb, 'h109be, 'h10bcb, 'h106fb, 'h1070b, 'h109bf, 'h1071b, 'h1072b, 'h109c0, 'h1073b, 'h1074b, 'h109c1, 'h1075b, 'h103bc, 'h1076b, 'h109c2, 'h1077b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078b, 'h109c3, 'h1079b, 'h10bcb, 'h107ab, 'h109c4, 'h107bb, 'h107cb, 'h109c5, 'h107db, 'h107eb, 'h109c6, 'h107fb, 'h1080b, 'h109c7, 'h103bc, 'h1081b, 'h1082b, 'h109c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083b, 'h1084b, 'h109c9, 'h10bcb, 'h1085b, 'h1086b, 'h109ca, 'h1087b, 'h1088b, 'h109cb, 'h1089b, 'h108ab, 'h109cc, 'h108bb, 'h103bc, 'h108cb, 'h109cd, 'h108db, 'h21f8e, 'h21f8f, 'h21f8d, 'h106eb, 'h109ce, 'h10bdb, 'h106fb, 'h1070b, 'h109cf, 'h1071b, 'h1072b, 'h109d0, 'h1073b, 'h1074b, 'h109d1, 'h1075b, 'h1076b, 'h109d2, 'h103bc, 'h1077b, 'h1078b, 'h109d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079b, 'h10bdb, 'h107ab, 'h109d4, 'h107bb, 'h107cb, 'h109d5, 'h107db, 'h107eb, 'h109d6, 'h107fb, 'h1080b, 'h109d7, 'h1081b, 'h103bc, 'h1082b, 'h109d8, 'h1083b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084b, 'h109d9, 'h10bdb, 'h1085b, 'h1086b, 'h109da, 'h1087b, 'h1088b, 'h109db, 'h1089b, 'h108ab, 'h109dc, 'h108bb, 'h108cb, 'h109dd, 'h103bc, 'h108db, 'h106eb, 'h109de, 'h10beb, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fb, 'h1070b, 'h109df, 'h1071b, 'h1072b, 'h109e0, 'h1073b, 'h1074b, 'h109e1, 'h1075b, 'h1076b, 'h109e2, 'h1077b, 'h103bc, 'h1078b, 'h109e3, 'h1079b, 'h10beb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ab, 'h109e4, 'h107bb, 'h107cb, 'h109e5, 'h107db, 'h107eb, 'h109e6, 'h107fb, 'h1080b, 'h109e7, 'h1081b, 'h1082b, 'h109e8, 'h103bc, 'h1083b, 'h1084b, 'h109e9, 'h10beb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085b, 'h1086b, 'h109ea, 'h1087b, 'h1088b, 'h109eb, 'h1089b, 'h108ab, 'h109ec, 'h108bb, 'h108cb, 'h109ed, 'h108db, 'h103bc, 'h106eb, 'h109ee, 'h10bfb, 'h106fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h109ef, 'h1071b, 'h1072b, 'h109f0, 'h1073b, 'h1074b, 'h109f1, 'h1075b, 'h1076b, 'h109f2, 'h1077b, 'h1078b, 'h109f3, 'h103bc, 'h1079b, 'h10bfb, 'h107ab, 'h109f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bb, 'h107cb, 'h109f5, 'h107db, 'h107eb, 'h109f6, 'h107fb, 'h1080b, 'h109f7, 'h1081b, 'h1082b, 'h109f8, 'h1083b, 'h103bc, 'h1084b, 'h109f9, 'h10bfb, 'h1085b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086b, 'h109fa, 'h1087b, 'h1088b, 'h109fb, 'h1089b, 'h108ab, 'h109fc, 'h108bb, 'h108cb, 'h109fd, 'h108db, 'h106eb, 'h109fe, 'h10c0b, 'h103bc, 'h106fb, 'h1070b, 'h109ff, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071b, 'h1072b, 'h10a00, 'h1073b, 'h1074b, 'h10a01, 'h1075b, 'h1076b, 'h10a02, 'h1077b, 'h1078b, 'h10a03, 'h1079b, 'h10c0b, 'h103bc, 'h107ab, 'h10a04, 'h107bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cb, 'h10a05, 'h107db, 'h107eb, 'h10a06, 'h107fb, 'h1080b, 'h10a07, 'h1081b, 'h1082b, 'h10a08, 'h1083b, 'h1084b, 'h10a09, 'h10c0b, 'h103bc, 'h1085b, 'h1086b, 'h10a0a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087b, 'h1088b, 'h10a0b, 'h1089b, 'h108ab, 'h10a0c, 'h108bb, 'h108cb, 'h10a0d, 'h108db, 'h106eb, 'h10a0e, 'h10c1b, 'h106fb, 'h103bc, 'h1070b, 'h10a0f, 'h1071b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072b, 'h10a10, 'h1073b, 'h1074b, 'h10a11, 'h1075b, 'h1076b, 'h10a12, 'h1077b, 'h1078b, 'h10a13, 'h1079b, 'h10c1b, 'h107ab, 'h10a14, 'h103bc, 'h107bb, 'h107cb, 'h10a15, 'h21f8e, 'h21f8f, 'h21f8d, 'h107db, 'h107eb, 'h10a16, 'h107fb, 'h1080b, 'h10a17, 'h1081b, 'h1082b, 'h10a18, 'h1083b, 'h1084b, 'h10a19, 'h10c1b, 'h1085b, 'h103bc, 'h1086b, 'h10a1a, 'h1087b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088b, 'h10a1b, 'h1089b, 'h108ab, 'h10a1c, 'h108bb, 'h108cb, 'h10a1d, 'h108db, 'h106eb, 'h10a1e, 'h10c2b, 'h106fb, 'h1070b, 'h10a1f, 'h103bc, 'h1071b, 'h1072b, 'h10a20, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h1074b, 'h10a21, 'h1075b, 'h1076b, 'h10a22, 'h1077b, 'h1078b, 'h10a23, 'h1079b, 'h10c2b, 'h107ab, 'h10a24, 'h107bb, 'h103bc, 'h107cb, 'h10a25, 'h107db, 'h21f8e, 'h21f8f, 'h21f8d, 'h107eb, 'h10a26, 'h107fb, 'h1080b, 'h10a27, 'h1081b, 'h1082b, 'h10a28, 'h1083b, 'h1084b, 'h10a29, 'h10c2b, 'h1085b, 'h1086b, 'h10a2a, 'h103bc, 'h1087b, 'h1088b, 'h10a2b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089b, 'h108ab, 'h10a2c, 'h108bb, 'h108cb, 'h10a2d, 'h108db, 'h106eb, 'h10a2e, 'h10c3b, 'h106fb, 'h1070b, 'h10a2f, 'h1071b, 'h103bc, 'h1072b, 'h10a30, 'h1073b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074b, 'h10a31, 'h1075b, 'h1076b, 'h10a32, 'h1077b, 'h1078b, 'h10a33, 'h1079b, 'h10c3b, 'h107ab, 'h10a34, 'h107bb, 'h107cb, 'h10a35, 'h103bc, 'h107db, 'h107eb, 'h10a36, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fb, 'h1080b, 'h10a37, 'h1081b, 'h1082b, 'h10a38, 'h1083b, 'h1084b, 'h10a39, 'h10c3b, 'h1085b, 'h1086b, 'h10a3a, 'h1087b, 'h103bc, 'h1088b, 'h10a3b, 'h1089b, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ab, 'h10a3c, 'h108bb, 'h108cb, 'h10a3d, 'h108db, 'h106eb, 'h10a3e, 'h10c4b, 'h106fb, 'h1070b, 'h10a3f, 'h1071b, 'h1072b, 'h10a40, 'h103bc, 'h1073b, 'h1074b, 'h10a41, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075b, 'h1076b, 'h10a42, 'h1077b, 'h1078b, 'h10a43, 'h1079b, 'h10c4b, 'h107ab, 'h10a44, 'h107bb, 'h107cb, 'h10a45, 'h107db, 'h103bc, 'h107eb, 'h10a46, 'h107fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080b, 'h10a47, 'h1081b, 'h1082b, 'h10a48, 'h1083b, 'h1084b, 'h10a49, 'h10c4b, 'h1085b, 'h1086b, 'h10a4a, 'h1087b, 'h1088b, 'h10a4b, 'h103bc, 'h1089b, 'h108ab, 'h10a4c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bb, 'h108cb, 'h10a4d, 'h108db, 'h106eb, 'h10a4e, 'h10c5b, 'h106fb, 'h1070b, 'h10a4f, 'h1071b, 'h1072b, 'h10a50, 'h1073b, 'h103bc, 'h1074b, 'h10a51, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076b, 'h10a52, 'h1077b, 'h1078b, 'h10a53, 'h1079b, 'h10c5b, 'h107ab, 'h10a54, 'h107bb, 'h107cb, 'h10a55, 'h107db, 'h107eb, 'h10a56, 'h103bc, 'h107fb, 'h1080b, 'h10a57, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081b, 'h1082b, 'h10a58, 'h1083b, 'h1084b, 'h10a59, 'h10c5b, 'h1085b, 'h1086b, 'h10a5a, 'h1087b, 'h1088b, 'h10a5b, 'h1089b, 'h103bc, 'h108ab, 'h10a5c, 'h108bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cb, 'h10a5d, 'h108db, 'h106eb, 'h10a5e, 'h10c6b, 'h106fb, 'h1070b, 'h10a5f, 'h1071b, 'h1072b, 'h10a60, 'h1073b, 'h1074b, 'h10a61, 'h103bc, 'h1075b, 'h1076b, 'h10a62, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077b, 'h1078b, 'h10a63, 'h1079b, 'h10c6b, 'h107ab, 'h10a64, 'h107bb, 'h107cb, 'h10a65, 'h107db, 'h107eb, 'h10a66, 'h107fb, 'h103bc, 'h1080b, 'h10a67, 'h1081b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082b, 'h10a68, 'h1083b, 'h1084b, 'h10a69, 'h10c6b, 'h1085b, 'h1086b, 'h10a6a, 'h1087b, 'h1088b, 'h10a6b, 'h1089b, 'h108ab, 'h10a6c, 'h103bc, 'h108bb, 'h108cb, 'h10a6d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108db, 'h106eb, 'h10a6e, 'h10c7b, 'h106fb, 'h1070b, 'h10a6f, 'h1071b, 'h1072b, 'h10a70, 'h1073b, 'h1074b, 'h10a71, 'h1075b, 'h103bc, 'h1076b, 'h10a72, 'h1077b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078b, 'h10a73, 'h1079b, 'h10c7b, 'h107ab, 'h10a74, 'h107bb, 'h107cb, 'h10a75, 'h107db, 'h107eb, 'h10a76, 'h107fb, 'h1080b, 'h10a77, 'h103bc, 'h1081b, 'h1082b, 'h10a78, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083b, 'h1084b, 'h10a79, 'h10c7b, 'h1085b, 'h1086b, 'h10a7a, 'h1087b, 'h1088b, 'h10a7b, 'h1089b, 'h108ab, 'h10a7c, 'h108bb, 'h103bc, 'h108cb, 'h10a7d, 'h108db, 'h21f8e, 'h21f8f, 'h21f8d, 'h106eb, 'h10a7e, 'h10c8b, 'h106fb, 'h1070b, 'h10a7f, 'h1071b, 'h1072b, 'h10a80, 'h1073b, 'h1074b, 'h10a81, 'h1075b, 'h1076b, 'h10a82, 'h103bc, 'h1077b, 'h1078b, 'h10a83, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079b, 'h10c8b, 'h107ab, 'h10a84, 'h107bb, 'h107cb, 'h10a85, 'h107db, 'h107eb, 'h10a86, 'h107fb, 'h1080b, 'h10a87, 'h1081b, 'h103bc, 'h1082b, 'h10a88, 'h1083b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084b, 'h10a89, 'h10c8b, 'h1085b, 'h1086b, 'h10a8a, 'h1087b, 'h1088b, 'h10a8b, 'h1089b, 'h108ab, 'h10a8c, 'h108bb, 'h108cb, 'h10a8d, 'h103bc, 'h108db, 'h106eb, 'h10a8e, 'h10c9b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fb, 'h1070b, 'h10a8f, 'h1071b, 'h1072b, 'h10a90, 'h1073b, 'h1074b, 'h10a91, 'h1075b, 'h1076b, 'h10a92, 'h1077b, 'h103bc, 'h1078b, 'h10a93, 'h1079b, 'h10c9b, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ab, 'h10a94, 'h107bb, 'h107cb, 'h10a95, 'h107db, 'h107eb, 'h10a96, 'h107fb, 'h1080b, 'h10a97, 'h1081b, 'h1082b, 'h10a98, 'h103bc, 'h1083b, 'h1084b, 'h10a99, 'h10c9b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085b, 'h1086b, 'h10a9a, 'h1087b, 'h1088b, 'h10a9b, 'h1089b, 'h108ab, 'h10a9c, 'h108bb, 'h108cb, 'h10a9d, 'h108db, 'h103bc, 'h106eb, 'h10a9e, 'h10cab, 'h106fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10a9f, 'h1071b, 'h1072b, 'h10aa0, 'h1073b, 'h1074b, 'h10aa1, 'h1075b, 'h1076b, 'h10aa2, 'h1077b, 'h1078b, 'h10aa3, 'h103bc, 'h1079b, 'h10cab, 'h107ab, 'h10aa4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bb, 'h107cb, 'h10aa5, 'h107db, 'h107eb, 'h10aa6, 'h107fb, 'h1080b, 'h10aa7, 'h1081b, 'h1082b, 'h10aa8, 'h1083b, 'h103bc, 'h1084b, 'h10aa9, 'h10cab, 'h1085b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086b, 'h10aaa, 'h1087b, 'h1088b, 'h10aab, 'h1089b, 'h108ab, 'h10aac, 'h108bb, 'h108cb, 'h10aad, 'h108db, 'h106eb, 'h10aae, 'h10cbb, 'h103bc, 'h106fb, 'h1070b, 'h10aaf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071b, 'h1072b, 'h10ab0, 'h1073b, 'h1074b, 'h10ab1, 'h1075b, 'h1076b, 'h10ab2, 'h1077b, 'h1078b, 'h10ab3, 'h1079b, 'h10cbb, 'h103bc, 'h107ab, 'h10ab4, 'h107bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cb, 'h10ab5, 'h107db, 'h107eb, 'h10ab6, 'h107fb, 'h1080b, 'h10ab7, 'h1081b, 'h1082b, 'h10ab8, 'h1083b, 'h1084b, 'h10ab9, 'h10cbb, 'h103bc, 'h1085b, 'h1086b, 'h10aba, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087b, 'h1088b, 'h10abb, 'h1089b, 'h108ab, 'h10abc, 'h108bb, 'h108cb, 'h10abd, 'h108db, 'h106eb, 'h10abe, 'h10ccb, 'h106fb, 'h103bc, 'h1070b, 'h10abf, 'h1071b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072b, 'h10ac0, 'h1073b, 'h1074b, 'h10ac1, 'h1075b, 'h1076b, 'h10ac2, 'h1077b, 'h1078b, 'h10ac3, 'h1079b, 'h10ccb, 'h107ab, 'h10ac4, 'h103bc, 'h107bb, 'h107cb, 'h10ac5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107db, 'h107eb, 'h10ac6, 'h107fb, 'h1080b, 'h10ac7, 'h1081b, 'h1082b, 'h10ac8, 'h1083b, 'h1084b, 'h10ac9, 'h10ccb, 'h1085b, 'h103bc, 'h1086b, 'h10aca, 'h1087b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088b, 'h10acb, 'h1089b, 'h108ab, 'h10acc, 'h108bb, 'h108cb, 'h10acd, 'h108db, 'h106eb, 'h10ace, 'h10cdb, 'h106fb, 'h1070b, 'h10acf, 'h103bc, 'h1071b, 'h1072b, 'h10ad0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h1074b, 'h10ad1, 'h1075b, 'h1076b, 'h10ad2, 'h1077b, 'h1078b, 'h10ad3, 'h1079b, 'h10cdb, 'h107ab, 'h10ad4, 'h107bb, 'h103bc, 'h107cb, 'h10ad5, 'h107db, 'h21f8e, 'h21f8f, 'h21f8d, 'h107eb, 'h10ad6, 'h107fb, 'h1080b, 'h10ad7, 'h1081b, 'h1082b, 'h10ad8, 'h1083b, 'h1084b, 'h10ad9, 'h10cdb, 'h1085b, 'h1086b, 'h10ada, 'h103bc, 'h1087b, 'h1088b, 'h10adb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089b, 'h108ab, 'h10adc, 'h108bb, 'h108cb, 'h10add, 'h108db, 'h106eb, 'h108de, 'h10aeb, 'h106fb, 'h1070b, 'h108df, 'h1071b, 'h103bc, 'h1072b, 'h108e0, 'h1073b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074b, 'h108e1, 'h1075b, 'h1076b, 'h108e2, 'h1077b, 'h1078b, 'h108e3, 'h1079b, 'h10aeb, 'h107ab, 'h108e4, 'h107bb, 'h107cb, 'h108e5, 'h103bc, 'h107db, 'h107eb, 'h108e6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fb, 'h1080b, 'h108e7, 'h1081b, 'h1082b, 'h108e8, 'h1083b, 'h1084b, 'h108e9, 'h10aeb, 'h1085b, 'h1086b, 'h108ea, 'h1087b, 'h103bc, 'h1088b, 'h108eb, 'h1089b, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ab, 'h108ec, 'h108bb, 'h108cb, 'h108ed, 'h108db, 'h106eb, 'h108ee, 'h10afb, 'h106fb, 'h1070b, 'h108ef, 'h1071b, 'h1072b, 'h108f0, 'h103bc, 'h1073b, 'h1074b, 'h108f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075b, 'h1076b, 'h108f2, 'h1077b, 'h1078b, 'h108f3, 'h1079b, 'h10afb, 'h107ab, 'h108f4, 'h107bb, 'h107cb, 'h108f5, 'h107db, 'h103bc, 'h107eb, 'h108f6, 'h107fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080b, 'h108f7, 'h1081b, 'h1082b, 'h108f8, 'h1083b, 'h1084b, 'h108f9, 'h10afb, 'h1085b, 'h1086b, 'h108fa, 'h1087b, 'h1088b, 'h108fb, 'h103bc, 'h1089b, 'h108ab, 'h108fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bb, 'h108cb, 'h108fd, 'h108db, 'h106eb, 'h108fe, 'h10b0b, 'h106fb, 'h1070b, 'h108ff, 'h1071b, 'h1072b, 'h10900, 'h1073b, 'h103bc, 'h1074b, 'h10901, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076b, 'h10902, 'h1077b, 'h1078b, 'h10903, 'h1079b, 'h10b0b, 'h107ab, 'h10904, 'h107bb, 'h107cb, 'h10905, 'h107db, 'h107eb, 'h10906, 'h103bc, 'h107fb, 'h1080b, 'h10907, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081b, 'h1082b, 'h10908, 'h1083b, 'h1084b, 'h10909, 'h10b0b, 'h1085b, 'h1086b, 'h1090a, 'h1087b, 'h1088b, 'h1090b, 'h1089b, 'h103bc, 'h108ab, 'h1090c, 'h108bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cb, 'h1090d, 'h108db, 'h106eb, 'h1090e, 'h10b1b, 'h106fb, 'h1070b, 'h1090f, 'h1071b, 'h1072b, 'h10910, 'h1073b, 'h1074b, 'h10911, 'h103bc, 'h1075b, 'h1076b, 'h10912, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077b, 'h1078b, 'h10913, 'h1079b, 'h10b1b, 'h107ab, 'h10914, 'h107bb, 'h107cb, 'h10915, 'h107db, 'h107eb, 'h10916, 'h107fb, 'h103bc, 'h1080b, 'h10917, 'h1081b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082b, 'h10918, 'h1083b, 'h1084b, 'h10919, 'h10b1b, 'h1085b, 'h1086b, 'h1091a, 'h1087b, 'h1088b, 'h1091b, 'h1089b, 'h108ab, 'h1091c, 'h103bc, 'h108bb, 'h108cb, 'h1091d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108db, 'h106eb, 'h1091e, 'h10b2b, 'h106fb, 'h1070b, 'h1091f, 'h1071b, 'h1072b, 'h10920, 'h1073b, 'h1074b, 'h10921, 'h1075b, 'h103bc, 'h1076b, 'h10922, 'h1077b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078b, 'h10923, 'h1079b, 'h10b2b, 'h107ab, 'h10924, 'h107bb, 'h107cb, 'h10925, 'h107db, 'h107eb, 'h10926, 'h107fb, 'h1080b, 'h10927, 'h103bc, 'h1081b, 'h1082b, 'h10928, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083b, 'h1084b, 'h10929, 'h10b2b, 'h1085b, 'h1086b, 'h1092a, 'h1087b, 'h1088b, 'h1092b, 'h1089b, 'h108ab, 'h1092c, 'h108bb, 'h103bc, 'h108cb, 'h1092d, 'h108db, 'h21f8e, 'h21f8f, 'h21f8d, 'h106eb, 'h1092e, 'h10b3b, 'h106fb, 'h1070b, 'h1092f, 'h1071b, 'h1072b, 'h10930, 'h1073b, 'h1074b, 'h10931, 'h1075b, 'h1076b, 'h10932, 'h103bc, 'h1077b, 'h1078b, 'h10933, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079b, 'h10b3b, 'h107ab, 'h10934, 'h107bb, 'h107cb, 'h10935, 'h107db, 'h107eb, 'h10936, 'h107fb, 'h1080b, 'h10937, 'h1081b, 'h103bc, 'h1082b, 'h10938, 'h1083b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084b, 'h10939, 'h10b3b, 'h1085b, 'h1086b, 'h1093a, 'h1087b, 'h1088b, 'h1093b, 'h1089b, 'h108ab, 'h1093c, 'h108bb, 'h108cb, 'h1093d, 'h103bc, 'h108db, 'h106eb, 'h1093e, 'h10b4b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fb, 'h1070b, 'h1093f, 'h1071b, 'h1072b, 'h10940, 'h1073b, 'h1074b, 'h10941, 'h1075b, 'h1076b, 'h10942, 'h1077b, 'h103bc, 'h1078b, 'h10943, 'h1079b, 'h10b4b, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ab, 'h10944, 'h107bb, 'h107cb, 'h10945, 'h107db, 'h107eb, 'h10946, 'h107fb, 'h1080b, 'h10947, 'h1081b, 'h1082b, 'h10948, 'h103bc, 'h1083b, 'h1084b, 'h10949, 'h10b4b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085b, 'h1086b, 'h1094a, 'h1087b, 'h1088b, 'h1094b, 'h1089b, 'h108ab, 'h1094c, 'h108bb, 'h108cb, 'h1094d, 'h108db, 'h103bc, 'h106eb, 'h1094e, 'h10b5b, 'h106fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h1094f, 'h1071b, 'h1072b, 'h10950, 'h1073b, 'h1074b, 'h10951, 'h1075b, 'h1076b, 'h10952, 'h1077b, 'h1078b, 'h10953, 'h103bc, 'h1079b, 'h10b5b, 'h107ab, 'h10954, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bb, 'h107cb, 'h10955, 'h107db, 'h107eb, 'h10956, 'h107fb, 'h1080b, 'h10957, 'h1081b, 'h1082b, 'h10958, 'h1083b, 'h103bc, 'h1084b, 'h10959, 'h10b5b, 'h1085b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086b, 'h1095a, 'h1087b, 'h1088b, 'h1095b, 'h1089b, 'h108ab, 'h1095c, 'h108bb, 'h108cb, 'h1095d, 'h108db, 'h106eb, 'h1095e, 'h10b6b, 'h103bc, 'h106fb, 'h1070b, 'h1095f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071b, 'h1072b, 'h10960, 'h1073b, 'h1074b, 'h10961, 'h1075b, 'h1076b, 'h10962, 'h1077b, 'h1078b, 'h10963, 'h1079b, 'h10b6b, 'h103bc, 'h107ab, 'h10964, 'h107bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cb, 'h10965, 'h107db, 'h107eb, 'h10966, 'h107fb, 'h1080b, 'h10967, 'h1081b, 'h1082b, 'h10968, 'h1083b, 'h1084b, 'h10969, 'h10b6b, 'h103bc, 'h1085b, 'h1086b, 'h1096a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087b, 'h1088b, 'h1096b, 'h1089b, 'h108ab, 'h1096c, 'h108bb, 'h108cb, 'h1096d, 'h108db, 'h106eb, 'h1096e, 'h10b7b, 'h106fb, 'h103bc, 'h1070b, 'h1096f, 'h1071b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072b, 'h10970, 'h1073b, 'h1074b, 'h10971, 'h1075b, 'h1076b, 'h10972, 'h1077b, 'h1078b, 'h10973, 'h1079b, 'h10b7b, 'h107ab, 'h10974, 'h103bc, 'h107bb, 'h107cb, 'h10975, 'h21f8e, 'h21f8f, 'h21f8d, 'h107db, 'h107eb, 'h10976, 'h107fb, 'h1080b, 'h10977, 'h1081b, 'h1082b, 'h10978, 'h1083b, 'h1084b, 'h10979, 'h10b7b, 'h1085b, 'h103bc, 'h1086b, 'h1097a, 'h1087b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088b, 'h1097b, 'h1089b, 'h108ab, 'h1097c, 'h108bb, 'h108cb, 'h1097d, 'h108db, 'h106eb, 'h1097e, 'h10b8b, 'h106fb, 'h1070b, 'h1097f, 'h103bc, 'h1071b, 'h1072b, 'h10980, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h1074b, 'h10981, 'h1075b, 'h1076b, 'h10982, 'h1077b, 'h1078b, 'h10983, 'h1079b, 'h10b8b, 'h107ab, 'h10984, 'h107bb, 'h103bc, 'h107cb, 'h10985, 'h107db, 'h21f8e, 'h21f8f, 'h21f8d, 'h107eb, 'h10986, 'h107fb, 'h1080b, 'h10987, 'h1081b, 'h1082b, 'h10988, 'h1083b, 'h1084b, 'h10989, 'h10b8b, 'h1085b, 'h1086b, 'h1098a, 'h103bc, 'h1087b, 'h1088b, 'h1098b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089b, 'h108ab, 'h1098c, 'h108bb, 'h108cb, 'h1098d, 'h108db, 'h106eb, 'h1098e, 'h10b9b, 'h106fb, 'h1070b, 'h1098f, 'h1071b, 'h103bc, 'h1072b, 'h10990, 'h1073b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074b, 'h10991, 'h1075b, 'h1076b, 'h10992, 'h1077b, 'h1078b, 'h10993, 'h1079b, 'h10b9b, 'h107ab, 'h10994, 'h107bb, 'h107cb, 'h10995, 'h103bc, 'h107db, 'h107eb, 'h10996, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fb, 'h1080b, 'h10997, 'h1081b, 'h1082b, 'h10998, 'h1083b, 'h1084b, 'h10999, 'h10b9b, 'h1085b, 'h1086b, 'h1099a, 'h1087b, 'h103bc, 'h1088b, 'h1099b, 'h1089b, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ab, 'h1099c, 'h108bb, 'h108cb, 'h1099d, 'h108db, 'h106eb, 'h1099e, 'h10bab, 'h106fb, 'h1070b, 'h1099f, 'h1071b, 'h1072b, 'h109a0, 'h103bc, 'h1073b, 'h1074b, 'h109a1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075b, 'h1076b, 'h109a2, 'h1077b, 'h1078b, 'h109a3, 'h1079b, 'h10bab, 'h107ab, 'h109a4, 'h107bb, 'h107cb, 'h109a5, 'h107db, 'h103bc, 'h107eb, 'h109a6, 'h107fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080b, 'h109a7, 'h1081b, 'h1082b, 'h109a8, 'h1083b, 'h1084b, 'h109a9, 'h10bab, 'h1085b, 'h1086b, 'h109aa, 'h1087b, 'h1088b, 'h109ab, 'h103bc, 'h1089b, 'h108ab, 'h109ac, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bb, 'h108cb, 'h109ad, 'h108db, 'h106eb, 'h109ae, 'h10bbb, 'h106fb, 'h1070b, 'h109af, 'h1071b, 'h1072b, 'h109b0, 'h1073b, 'h103bc, 'h1074b, 'h109b1, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076b, 'h109b2, 'h1077b, 'h1078b, 'h109b3, 'h1079b, 'h10bbb, 'h107ab, 'h109b4, 'h107bb, 'h107cb, 'h109b5, 'h107db, 'h107eb, 'h109b6, 'h103bc, 'h107fb, 'h1080b, 'h109b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081b, 'h1082b, 'h109b8, 'h1083b, 'h1084b, 'h109b9, 'h10bbb, 'h1085b, 'h1086b, 'h109ba, 'h1087b, 'h1088b, 'h109bb, 'h1089b, 'h103bc, 'h108ab, 'h109bc, 'h108bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cb, 'h109bd, 'h108db, 'h106eb, 'h109be, 'h10bcb, 'h106fb, 'h1070b, 'h109bf, 'h1071b, 'h1072b, 'h109c0, 'h1073b, 'h1074b, 'h109c1, 'h103bc, 'h1075b, 'h1076b, 'h109c2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077b, 'h1078b, 'h109c3, 'h1079b, 'h10bcb, 'h107ab, 'h109c4, 'h107bb, 'h107cb, 'h109c5, 'h107db, 'h107eb, 'h109c6, 'h107fb, 'h103bc, 'h1080b, 'h109c7, 'h1081b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082b, 'h109c8, 'h1083b, 'h1084b, 'h109c9, 'h10bcb, 'h1085b, 'h1086b, 'h109ca, 'h1087b, 'h1088b, 'h109cb, 'h1089b, 'h108ab, 'h109cc, 'h103bc, 'h108bb, 'h108cb, 'h109cd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108db, 'h106eb, 'h109ce, 'h10bdb, 'h106fb, 'h1070b, 'h109cf, 'h1071b, 'h1072b, 'h109d0, 'h1073b, 'h1074b, 'h109d1, 'h1075b, 'h103bc, 'h1076b, 'h109d2, 'h1077b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078b, 'h109d3, 'h1079b, 'h10bdb, 'h107ab, 'h109d4, 'h107bb, 'h107cb, 'h109d5, 'h107db, 'h107eb, 'h109d6, 'h107fb, 'h1080b, 'h109d7, 'h103bc, 'h1081b, 'h1082b, 'h109d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083b, 'h1084b, 'h109d9, 'h10bdb, 'h1085b, 'h1086b, 'h109da, 'h1087b, 'h1088b, 'h109db, 'h1089b, 'h108ab, 'h109dc, 'h108bb, 'h103bc, 'h108cb, 'h109dd, 'h108db, 'h21f8e, 'h21f8f, 'h21f8d, 'h106eb, 'h109de, 'h10beb, 'h106fb, 'h1070b, 'h109df, 'h1071b, 'h1072b, 'h109e0, 'h1073b, 'h1074b, 'h109e1, 'h1075b, 'h1076b, 'h109e2, 'h103bc, 'h1077b, 'h1078b, 'h109e3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079b, 'h10beb, 'h107ab, 'h109e4, 'h107bb, 'h107cb, 'h109e5, 'h107db, 'h107eb, 'h109e6, 'h107fb, 'h1080b, 'h109e7, 'h1081b, 'h103bc, 'h1082b, 'h109e8, 'h1083b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084b, 'h109e9, 'h10beb, 'h1085b, 'h1086b, 'h109ea, 'h1087b, 'h1088b, 'h109eb, 'h1089b, 'h108ab, 'h109ec, 'h108bb, 'h108cb, 'h109ed, 'h103bc, 'h108db, 'h106eb, 'h109ee, 'h10bfb, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fb, 'h1070b, 'h109ef, 'h1071b, 'h1072b, 'h109f0, 'h1073b, 'h1074b, 'h109f1, 'h1075b, 'h1076b, 'h109f2, 'h1077b, 'h103bc, 'h1078b, 'h109f3, 'h1079b, 'h10bfb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ab, 'h109f4, 'h107bb, 'h107cb, 'h109f5, 'h107db, 'h107eb, 'h109f6, 'h107fb, 'h1080b, 'h109f7, 'h1081b, 'h1082b, 'h109f8, 'h103bc, 'h1083b, 'h1084b, 'h109f9, 'h10bfb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085b, 'h1086b, 'h109fa, 'h1087b, 'h1088b, 'h109fb, 'h1089b, 'h108ab, 'h109fc, 'h108bb, 'h108cb, 'h109fd, 'h108db, 'h103bc, 'h106eb, 'h109fe, 'h10c0b, 'h106fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h109ff, 'h1071b, 'h1072b, 'h10a00, 'h1073b, 'h1074b, 'h10a01, 'h1075b, 'h1076b, 'h10a02, 'h1077b, 'h1078b, 'h10a03, 'h103bc, 'h1079b, 'h10c0b, 'h107ab, 'h10a04, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bb, 'h107cb, 'h10a05, 'h107db, 'h107eb, 'h10a06, 'h107fb, 'h1080b, 'h10a07, 'h1081b, 'h1082b, 'h10a08, 'h1083b, 'h103bc, 'h1084b, 'h10a09, 'h10c0b, 'h1085b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086b, 'h10a0a, 'h1087b, 'h1088b, 'h10a0b, 'h1089b, 'h108ab, 'h10a0c, 'h108bb, 'h108cb, 'h10a0d, 'h108db, 'h106eb, 'h10a0e, 'h10c1b, 'h103bc, 'h106fb, 'h1070b, 'h10a0f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071b, 'h1072b, 'h10a10, 'h1073b, 'h1074b, 'h10a11, 'h1075b, 'h1076b, 'h10a12, 'h1077b, 'h1078b, 'h10a13, 'h1079b, 'h10c1b, 'h103bc, 'h107ab, 'h10a14, 'h107bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cb, 'h10a15, 'h107db, 'h107eb, 'h10a16, 'h107fb, 'h1080b, 'h10a17, 'h1081b, 'h1082b, 'h10a18, 'h1083b, 'h1084b, 'h10a19, 'h10c1b, 'h103bc, 'h1085b, 'h1086b, 'h10a1a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087b, 'h1088b, 'h10a1b, 'h1089b, 'h108ab, 'h10a1c, 'h108bb, 'h108cb, 'h10a1d, 'h108db, 'h106eb, 'h10a1e, 'h10c2b, 'h106fb, 'h103bc, 'h1070b, 'h10a1f, 'h1071b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072b, 'h10a20, 'h1073b, 'h1074b, 'h10a21, 'h1075b, 'h1076b, 'h10a22, 'h1077b, 'h1078b, 'h10a23, 'h1079b, 'h10c2b, 'h107ab, 'h10a24, 'h103bc, 'h107bb, 'h107cb, 'h10a25, 'h21f8e, 'h21f8f, 'h21f8d, 'h107db, 'h107eb, 'h10a26, 'h107fb, 'h1080b, 'h10a27, 'h1081b, 'h1082b, 'h10a28, 'h1083b, 'h1084b, 'h10a29, 'h10c2b, 'h1085b, 'h103bc, 'h1086b, 'h10a2a, 'h1087b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088b, 'h10a2b, 'h1089b, 'h108ab, 'h10a2c, 'h108bb, 'h108cb, 'h10a2d, 'h108db, 'h106eb, 'h10a2e, 'h10c3b, 'h106fb, 'h1070b, 'h10a2f, 'h103bc, 'h1071b, 'h1072b, 'h10a30, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h1074b, 'h10a31, 'h1075b, 'h1076b, 'h10a32, 'h1077b, 'h1078b, 'h10a33, 'h1079b, 'h10c3b, 'h107ab, 'h10a34, 'h107bb, 'h103bc, 'h107cb, 'h10a35, 'h107db, 'h21f8e, 'h21f8f, 'h21f8d, 'h107eb, 'h10a36, 'h107fb, 'h1080b, 'h10a37, 'h1081b, 'h1082b, 'h10a38, 'h1083b, 'h1084b, 'h10a39, 'h10c3b, 'h1085b, 'h1086b, 'h10a3a, 'h103bc, 'h1087b, 'h1088b, 'h10a3b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089b, 'h108ab, 'h10a3c, 'h108bb, 'h108cb, 'h10a3d, 'h108db, 'h106eb, 'h10a3e, 'h10c4b, 'h106fb, 'h1070b, 'h10a3f, 'h1071b, 'h103bc, 'h1072b, 'h10a40, 'h1073b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074b, 'h10a41, 'h1075b, 'h1076b, 'h10a42, 'h1077b, 'h1078b, 'h10a43, 'h1079b, 'h10c4b, 'h107ab, 'h10a44, 'h107bb, 'h107cb, 'h10a45, 'h103bc, 'h107db, 'h107eb, 'h10a46, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fb, 'h1080b, 'h10a47, 'h1081b, 'h1082b, 'h10a48, 'h1083b, 'h1084b, 'h10a49, 'h10c4b, 'h1085b, 'h1086b, 'h10a4a, 'h1087b, 'h103bc, 'h1088b, 'h10a4b, 'h1089b, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ab, 'h10a4c, 'h108bb, 'h108cb, 'h10a4d, 'h108db, 'h106eb, 'h10a4e, 'h10c5b, 'h106fb, 'h1070b, 'h10a4f, 'h1071b, 'h1072b, 'h10a50, 'h103bc, 'h1073b, 'h1074b, 'h10a51, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075b, 'h1076b, 'h10a52, 'h1077b, 'h1078b, 'h10a53, 'h1079b, 'h10c5b, 'h107ab, 'h10a54, 'h107bb, 'h107cb, 'h10a55, 'h107db, 'h103bc, 'h107eb, 'h10a56, 'h107fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080b, 'h10a57, 'h1081b, 'h1082b, 'h10a58, 'h1083b, 'h1084b, 'h10a59, 'h10c5b, 'h1085b, 'h1086b, 'h10a5a, 'h1087b, 'h1088b, 'h10a5b, 'h103bc, 'h1089b, 'h108ab, 'h10a5c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bb, 'h108cb, 'h10a5d, 'h108db, 'h106eb, 'h10a5e, 'h10c6b, 'h106fb, 'h1070b, 'h10a5f, 'h1071b, 'h1072b, 'h10a60, 'h1073b, 'h103bc, 'h1074b, 'h10a61, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076b, 'h10a62, 'h1077b, 'h1078b, 'h10a63, 'h1079b, 'h10c6b, 'h107ab, 'h10a64, 'h107bb, 'h107cb, 'h10a65, 'h107db, 'h107eb, 'h10a66, 'h103bc, 'h107fb, 'h1080b, 'h10a67, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081b, 'h1082b, 'h10a68, 'h1083b, 'h1084b, 'h10a69, 'h10c6b, 'h1085b, 'h1086b, 'h10a6a, 'h1087b, 'h1088b, 'h10a6b, 'h1089b, 'h103bc, 'h108ab, 'h10a6c, 'h108bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cb, 'h10a6d, 'h108db, 'h106eb, 'h10a6e, 'h10c7b, 'h106fb, 'h1070b, 'h10a6f, 'h1071b, 'h1072b, 'h10a70, 'h1073b, 'h1074b, 'h10a71, 'h103bc, 'h1075b, 'h1076b, 'h10a72, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077b, 'h1078b, 'h10a73, 'h1079b, 'h10c7b, 'h107ab, 'h10a74, 'h107bb, 'h107cb, 'h10a75, 'h107db, 'h107eb, 'h10a76, 'h107fb, 'h103bc, 'h1080b, 'h10a77, 'h1081b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082b, 'h10a78, 'h1083b, 'h1084b, 'h10a79, 'h10c7b, 'h1085b, 'h1086b, 'h10a7a, 'h1087b, 'h1088b, 'h10a7b, 'h1089b, 'h108ab, 'h10a7c, 'h103bc, 'h108bb, 'h108cb, 'h10a7d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108db, 'h106eb, 'h10a7e, 'h10c8b, 'h106fb, 'h1070b, 'h10a7f, 'h1071b, 'h1072b, 'h10a80, 'h1073b, 'h1074b, 'h10a81, 'h1075b, 'h103bc, 'h1076b, 'h10a82, 'h1077b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078b, 'h10a83, 'h1079b, 'h10c8b, 'h107ab, 'h10a84, 'h107bb, 'h107cb, 'h10a85, 'h107db, 'h107eb, 'h10a86, 'h107fb, 'h1080b, 'h10a87, 'h103bc, 'h1081b, 'h1082b, 'h10a88, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083b, 'h1084b, 'h10a89, 'h10c8b, 'h1085b, 'h1086b, 'h10a8a, 'h1087b, 'h1088b, 'h10a8b, 'h1089b, 'h108ab, 'h10a8c, 'h108bb, 'h103bc, 'h108cb, 'h10a8d, 'h108db, 'h21f8e, 'h21f8f, 'h21f8d, 'h106eb, 'h10a8e, 'h10c9b, 'h106fb, 'h1070b, 'h10a8f, 'h1071b, 'h1072b, 'h10a90, 'h1073b, 'h1074b, 'h10a91, 'h1075b, 'h1076b, 'h10a92, 'h103bc, 'h1077b, 'h1078b, 'h10a93, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079b, 'h10c9b, 'h107ab, 'h10a94, 'h107bb, 'h107cb, 'h10a95, 'h107db, 'h107eb, 'h10a96, 'h107fb, 'h1080b, 'h10a97, 'h1081b, 'h103bc, 'h1082b, 'h10a98, 'h1083b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084b, 'h10a99, 'h10c9b, 'h1085b, 'h1086b, 'h10a9a, 'h1087b, 'h1088b, 'h10a9b, 'h1089b, 'h108ab, 'h10a9c, 'h108bb, 'h108cb, 'h10a9d, 'h103bc, 'h108db, 'h106eb, 'h10a9e, 'h10cab, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fb, 'h1070b, 'h10a9f, 'h1071b, 'h1072b, 'h10aa0, 'h1073b, 'h1074b, 'h10aa1, 'h1075b, 'h1076b, 'h10aa2, 'h1077b, 'h103bc, 'h1078b, 'h10aa3, 'h1079b, 'h10cab, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ab, 'h10aa4, 'h107bb, 'h107cb, 'h10aa5, 'h107db, 'h107eb, 'h10aa6, 'h107fb, 'h1080b, 'h10aa7, 'h1081b, 'h1082b, 'h10aa8, 'h103bc, 'h1083b, 'h1084b, 'h10aa9, 'h10cab, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085b, 'h1086b, 'h10aaa, 'h1087b, 'h1088b, 'h10aab, 'h1089b, 'h108ab, 'h10aac, 'h108bb, 'h108cb, 'h10aad, 'h108db, 'h103bc, 'h106eb, 'h10aae, 'h10cbb, 'h106fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10aaf, 'h1071b, 'h1072b, 'h10ab0, 'h1073b, 'h1074b, 'h10ab1, 'h1075b, 'h1076b, 'h10ab2, 'h1077b, 'h1078b, 'h10ab3, 'h103bc, 'h1079b, 'h10cbb, 'h107ab, 'h10ab4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bb, 'h107cb, 'h10ab5, 'h107db, 'h107eb, 'h10ab6, 'h107fb, 'h1080b, 'h10ab7, 'h1081b, 'h1082b, 'h10ab8, 'h1083b, 'h103bc, 'h1084b, 'h10ab9, 'h10cbb, 'h1085b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086b, 'h10aba, 'h1087b, 'h1088b, 'h10abb, 'h1089b, 'h108ab, 'h10abc, 'h108bb, 'h108cb, 'h10abd, 'h108db, 'h106eb, 'h10abe, 'h10ccb, 'h103bc, 'h106fb, 'h1070b, 'h10abf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071b, 'h1072b, 'h10ac0, 'h1073b, 'h1074b, 'h10ac1, 'h1075b, 'h1076b, 'h10ac2, 'h1077b, 'h1078b, 'h10ac3, 'h1079b, 'h10ccb, 'h103bc, 'h107ab, 'h10ac4, 'h107bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cb, 'h10ac5, 'h107db, 'h107eb, 'h10ac6, 'h107fb, 'h1080b, 'h10ac7, 'h1081b, 'h1082b, 'h10ac8, 'h1083b, 'h1084b, 'h10ac9, 'h10ccb, 'h103bc, 'h1085b, 'h1086b, 'h10aca, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087b, 'h1088b, 'h10acb, 'h1089b, 'h108ab, 'h10acc, 'h108bb, 'h108cb, 'h10acd, 'h108db, 'h106eb, 'h10ace, 'h10cdb, 'h106fb, 'h103bc, 'h1070b, 'h10acf, 'h1071b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072b, 'h10ad0, 'h1073b, 'h1074b, 'h10ad1, 'h1075b, 'h1076b, 'h10ad2, 'h1077b, 'h1078b, 'h10ad3, 'h1079b, 'h10cdb, 'h107ab, 'h10ad4, 'h103bc, 'h107bb, 'h107cb, 'h10ad5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107db, 'h107eb, 'h10ad6, 'h107fb, 'h1080b, 'h10ad7, 'h1081b, 'h1082b, 'h10ad8, 'h1083b, 'h1084b, 'h10ad9, 'h10cdb, 'h1085b, 'h103bc, 'h1086b, 'h10ada, 'h1087b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088b, 'h10adb, 'h1089b, 'h108ab, 'h10adc, 'h108bb, 'h108cb, 'h10add, 'h108db, 'h106ec, 'h108de, 'h10aec, 'h106fc, 'h1070c, 'h108df, 'h103bc, 'h1071c, 'h1072c, 'h108e0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h1074c, 'h108e1, 'h1075c, 'h1076c, 'h108e2, 'h1077c, 'h1078c, 'h108e3, 'h1079c, 'h10aec, 'h107ac, 'h108e4, 'h107bc, 'h103bc, 'h107cc, 'h108e5, 'h107dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ec, 'h108e6, 'h107fc, 'h1080c, 'h108e7, 'h1081c, 'h1082c, 'h108e8, 'h1083c, 'h1084c, 'h108e9, 'h10aec, 'h1085c, 'h1086c, 'h108ea, 'h103bc, 'h1087c, 'h1088c, 'h108eb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089c, 'h108ac, 'h108ec, 'h108bc, 'h108cc, 'h108ed, 'h108dc, 'h106ec, 'h108ee, 'h10afc, 'h106fc, 'h1070c, 'h108ef, 'h1071c, 'h103bc, 'h1072c, 'h108f0, 'h1073c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074c, 'h108f1, 'h1075c, 'h1076c, 'h108f2, 'h1077c, 'h1078c, 'h108f3, 'h1079c, 'h10afc, 'h107ac, 'h108f4, 'h107bc, 'h107cc, 'h108f5, 'h103bc, 'h107dc, 'h107ec, 'h108f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fc, 'h1080c, 'h108f7, 'h1081c, 'h1082c, 'h108f8, 'h1083c, 'h1084c, 'h108f9, 'h10afc, 'h1085c, 'h1086c, 'h108fa, 'h1087c, 'h103bc, 'h1088c, 'h108fb, 'h1089c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ac, 'h108fc, 'h108bc, 'h108cc, 'h108fd, 'h108dc, 'h106ec, 'h108fe, 'h10b0c, 'h106fc, 'h1070c, 'h108ff, 'h1071c, 'h1072c, 'h10900, 'h103bc, 'h1073c, 'h1074c, 'h10901, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075c, 'h1076c, 'h10902, 'h1077c, 'h1078c, 'h10903, 'h1079c, 'h10b0c, 'h107ac, 'h10904, 'h107bc, 'h107cc, 'h10905, 'h107dc, 'h103bc, 'h107ec, 'h10906, 'h107fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080c, 'h10907, 'h1081c, 'h1082c, 'h10908, 'h1083c, 'h1084c, 'h10909, 'h10b0c, 'h1085c, 'h1086c, 'h1090a, 'h1087c, 'h1088c, 'h1090b, 'h103bc, 'h1089c, 'h108ac, 'h1090c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bc, 'h108cc, 'h1090d, 'h108dc, 'h106ec, 'h1090e, 'h10b1c, 'h106fc, 'h1070c, 'h1090f, 'h1071c, 'h1072c, 'h10910, 'h1073c, 'h103bc, 'h1074c, 'h10911, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076c, 'h10912, 'h1077c, 'h1078c, 'h10913, 'h1079c, 'h10b1c, 'h107ac, 'h10914, 'h107bc, 'h107cc, 'h10915, 'h107dc, 'h107ec, 'h10916, 'h103bc, 'h107fc, 'h1080c, 'h10917, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081c, 'h1082c, 'h10918, 'h1083c, 'h1084c, 'h10919, 'h10b1c, 'h1085c, 'h1086c, 'h1091a, 'h1087c, 'h1088c, 'h1091b, 'h1089c, 'h103bc, 'h108ac, 'h1091c, 'h108bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cc, 'h1091d, 'h108dc, 'h106ec, 'h1091e, 'h10b2c, 'h106fc, 'h1070c, 'h1091f, 'h1071c, 'h1072c, 'h10920, 'h1073c, 'h1074c, 'h10921, 'h103bc, 'h1075c, 'h1076c, 'h10922, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077c, 'h1078c, 'h10923, 'h1079c, 'h10b2c, 'h107ac, 'h10924, 'h107bc, 'h107cc, 'h10925, 'h107dc, 'h107ec, 'h10926, 'h107fc, 'h103bc, 'h1080c, 'h10927, 'h1081c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082c, 'h10928, 'h1083c, 'h1084c, 'h10929, 'h10b2c, 'h1085c, 'h1086c, 'h1092a, 'h1087c, 'h1088c, 'h1092b, 'h1089c, 'h108ac, 'h1092c, 'h103bc, 'h108bc, 'h108cc, 'h1092d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108dc, 'h106ec, 'h1092e, 'h10b3c, 'h106fc, 'h1070c, 'h1092f, 'h1071c, 'h1072c, 'h10930, 'h1073c, 'h1074c, 'h10931, 'h1075c, 'h103bc, 'h1076c, 'h10932, 'h1077c, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078c, 'h10933, 'h1079c, 'h10b3c, 'h107ac, 'h10934, 'h107bc, 'h107cc, 'h10935, 'h107dc, 'h107ec, 'h10936, 'h107fc, 'h1080c, 'h10937, 'h103bc, 'h1081c, 'h1082c, 'h10938, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083c, 'h1084c, 'h10939, 'h10b3c, 'h1085c, 'h1086c, 'h1093a, 'h1087c, 'h1088c, 'h1093b, 'h1089c, 'h108ac, 'h1093c, 'h108bc, 'h103bc, 'h108cc, 'h1093d, 'h108dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ec, 'h1093e, 'h10b4c, 'h106fc, 'h1070c, 'h1093f, 'h1071c, 'h1072c, 'h10940, 'h1073c, 'h1074c, 'h10941, 'h1075c, 'h1076c, 'h10942, 'h103bc, 'h1077c, 'h1078c, 'h10943, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079c};
	int DATA7 [7*SIZE-1:0] = {DATA6, DATA0};
	
endpackage
