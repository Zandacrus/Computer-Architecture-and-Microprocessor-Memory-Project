

package MATRIX_MULTIPLY_32_PKG_6;
	
	import MATRIX_MULTIPLY_32_PKG_5::DATA5;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h106e7, 'h10a4e, 'h10c57, 'h106f7, 'h103bc, 'h10707, 'h10a4f, 'h10717, 'h21f8e, 'h21f8f, 'h21f8d, 'h10727, 'h10a50, 'h10737, 'h10747, 'h10a51, 'h10757, 'h10767, 'h10a52, 'h10777, 'h10787, 'h10a53, 'h10797, 'h10c57, 'h107a7, 'h10a54, 'h103bc, 'h107b7, 'h107c7, 'h10a55, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d7, 'h107e7, 'h10a56, 'h107f7, 'h10807, 'h10a57, 'h10817, 'h10827, 'h10a58, 'h10837, 'h10847, 'h10a59, 'h10c57, 'h10857, 'h103bc, 'h10867, 'h10a5a, 'h10877, 'h21f8e, 'h21f8f, 'h21f8d, 'h10887, 'h10a5b, 'h10897, 'h108a7, 'h10a5c, 'h108b7, 'h108c7, 'h10a5d, 'h108d7, 'h106e7, 'h10a5e, 'h10c67, 'h106f7, 'h10707, 'h10a5f, 'h103bc, 'h10717, 'h10727, 'h10a60, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h10747, 'h10a61, 'h10757, 'h10767, 'h10a62, 'h10777, 'h10787, 'h10a63, 'h10797, 'h10c67, 'h107a7, 'h10a64, 'h107b7, 'h103bc, 'h107c7, 'h10a65, 'h107d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e7, 'h10a66, 'h107f7, 'h10807, 'h10a67, 'h10817, 'h10827, 'h10a68, 'h10837, 'h10847, 'h10a69, 'h10c67, 'h10857, 'h10867, 'h10a6a, 'h103bc, 'h10877, 'h10887, 'h10a6b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10897, 'h108a7, 'h10a6c, 'h108b7, 'h108c7, 'h10a6d, 'h108d7, 'h106e7, 'h10a6e, 'h10c77, 'h106f7, 'h10707, 'h10a6f, 'h10717, 'h103bc, 'h10727, 'h10a70, 'h10737, 'h21f8e, 'h21f8f, 'h21f8d, 'h10747, 'h10a71, 'h10757, 'h10767, 'h10a72, 'h10777, 'h10787, 'h10a73, 'h10797, 'h10c77, 'h107a7, 'h10a74, 'h107b7, 'h107c7, 'h10a75, 'h103bc, 'h107d7, 'h107e7, 'h10a76, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f7, 'h10807, 'h10a77, 'h10817, 'h10827, 'h10a78, 'h10837, 'h10847, 'h10a79, 'h10c77, 'h10857, 'h10867, 'h10a7a, 'h10877, 'h103bc, 'h10887, 'h10a7b, 'h10897, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a7, 'h10a7c, 'h108b7, 'h108c7, 'h10a7d, 'h108d7, 'h106e7, 'h10a7e, 'h10c87, 'h106f7, 'h10707, 'h10a7f, 'h10717, 'h10727, 'h10a80, 'h103bc, 'h10737, 'h10747, 'h10a81, 'h21f8e, 'h21f8f, 'h21f8d, 'h10757, 'h10767, 'h10a82, 'h10777, 'h10787, 'h10a83, 'h10797, 'h10c87, 'h107a7, 'h10a84, 'h107b7, 'h107c7, 'h10a85, 'h107d7, 'h103bc, 'h107e7, 'h10a86, 'h107f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10807, 'h10a87, 'h10817, 'h10827, 'h10a88, 'h10837, 'h10847, 'h10a89, 'h10c87, 'h10857, 'h10867, 'h10a8a, 'h10877, 'h10887, 'h10a8b, 'h103bc, 'h10897, 'h108a7, 'h10a8c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b7, 'h108c7, 'h10a8d, 'h108d7, 'h106e7, 'h10a8e, 'h10c97, 'h106f7, 'h10707, 'h10a8f, 'h10717, 'h10727, 'h10a90, 'h10737, 'h103bc, 'h10747, 'h10a91, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h10767, 'h10a92, 'h10777, 'h10787, 'h10a93, 'h10797, 'h10c97, 'h107a7, 'h10a94, 'h107b7, 'h107c7, 'h10a95, 'h107d7, 'h107e7, 'h10a96, 'h103bc, 'h107f7, 'h10807, 'h10a97, 'h21f8e, 'h21f8f, 'h21f8d, 'h10817, 'h10827, 'h10a98, 'h10837, 'h10847, 'h10a99, 'h10c97, 'h10857, 'h10867, 'h10a9a, 'h10877, 'h10887, 'h10a9b, 'h10897, 'h103bc, 'h108a7, 'h10a9c, 'h108b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c7, 'h10a9d, 'h108d7, 'h106e7, 'h10a9e, 'h10ca7, 'h106f7, 'h10707, 'h10a9f, 'h10717, 'h10727, 'h10aa0, 'h10737, 'h10747, 'h10aa1, 'h103bc, 'h10757, 'h10767, 'h10aa2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10777, 'h10787, 'h10aa3, 'h10797, 'h10ca7, 'h107a7, 'h10aa4, 'h107b7, 'h107c7, 'h10aa5, 'h107d7, 'h107e7, 'h10aa6, 'h107f7, 'h103bc, 'h10807, 'h10aa7, 'h10817, 'h21f8e, 'h21f8f, 'h21f8d, 'h10827, 'h10aa8, 'h10837, 'h10847, 'h10aa9, 'h10ca7, 'h10857, 'h10867, 'h10aaa, 'h10877, 'h10887, 'h10aab, 'h10897, 'h108a7, 'h10aac, 'h103bc, 'h108b7, 'h108c7, 'h10aad, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d7, 'h106e7, 'h10aae, 'h10cb7, 'h106f7, 'h10707, 'h10aaf, 'h10717, 'h10727, 'h10ab0, 'h10737, 'h10747, 'h10ab1, 'h10757, 'h103bc, 'h10767, 'h10ab2, 'h10777, 'h21f8e, 'h21f8f, 'h21f8d, 'h10787, 'h10ab3, 'h10797, 'h10cb7, 'h107a7, 'h10ab4, 'h107b7, 'h107c7, 'h10ab5, 'h107d7, 'h107e7, 'h10ab6, 'h107f7, 'h10807, 'h10ab7, 'h103bc, 'h10817, 'h10827, 'h10ab8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10837, 'h10847, 'h10ab9, 'h10cb7, 'h10857, 'h10867, 'h10aba, 'h10877, 'h10887, 'h10abb, 'h10897, 'h108a7, 'h10abc, 'h108b7, 'h103bc, 'h108c7, 'h10abd, 'h108d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e7, 'h10abe, 'h10cc7, 'h106f7, 'h10707, 'h10abf, 'h10717, 'h10727, 'h10ac0, 'h10737, 'h10747, 'h10ac1, 'h10757, 'h10767, 'h10ac2, 'h103bc, 'h10777, 'h10787, 'h10ac3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10797, 'h10cc7, 'h107a7, 'h10ac4, 'h107b7, 'h107c7, 'h10ac5, 'h107d7, 'h107e7, 'h10ac6, 'h107f7, 'h10807, 'h10ac7, 'h10817, 'h103bc, 'h10827, 'h10ac8, 'h10837, 'h21f8e, 'h21f8f, 'h21f8d, 'h10847, 'h10ac9, 'h10cc7, 'h10857, 'h10867, 'h10aca, 'h10877, 'h10887, 'h10acb, 'h10897, 'h108a7, 'h10acc, 'h108b7, 'h108c7, 'h10acd, 'h103bc, 'h108d7, 'h106e7, 'h10ace, 'h10cd7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f7, 'h10707, 'h10acf, 'h10717, 'h10727, 'h10ad0, 'h10737, 'h10747, 'h10ad1, 'h10757, 'h10767, 'h10ad2, 'h10777, 'h103bc, 'h10787, 'h10ad3, 'h10797, 'h10cd7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a7, 'h10ad4, 'h107b7, 'h107c7, 'h10ad5, 'h107d7, 'h107e7, 'h10ad6, 'h107f7, 'h10807, 'h10ad7, 'h10817, 'h10827, 'h10ad8, 'h103bc, 'h10837, 'h10847, 'h10ad9, 'h10cd7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10857, 'h10867, 'h10ada, 'h10877, 'h10887, 'h10adb, 'h10897, 'h108a7, 'h10adc, 'h108b7, 'h108c7, 'h10add, 'h108d7, 'h103bc, 'h106e8, 'h108de, 'h10ae8, 'h106f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h108df, 'h10718, 'h10728, 'h108e0, 'h10738, 'h10748, 'h108e1, 'h10758, 'h10768, 'h108e2, 'h10778, 'h10788, 'h108e3, 'h103bc, 'h10798, 'h10ae8, 'h107a8, 'h108e4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b8, 'h107c8, 'h108e5, 'h107d8, 'h107e8, 'h108e6, 'h107f8, 'h10808, 'h108e7, 'h10818, 'h10828, 'h108e8, 'h10838, 'h103bc, 'h10848, 'h108e9, 'h10ae8, 'h10858, 'h21f8e, 'h21f8f, 'h21f8d, 'h10868, 'h108ea, 'h10878, 'h10888, 'h108eb, 'h10898, 'h108a8, 'h108ec, 'h108b8, 'h108c8, 'h108ed, 'h108d8, 'h106e8, 'h108ee, 'h10af8, 'h103bc, 'h106f8, 'h10708, 'h108ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h10718, 'h10728, 'h108f0, 'h10738, 'h10748, 'h108f1, 'h10758, 'h10768, 'h108f2, 'h10778, 'h10788, 'h108f3, 'h10798, 'h10af8, 'h103bc, 'h107a8, 'h108f4, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c8, 'h108f5, 'h107d8, 'h107e8, 'h108f6, 'h107f8, 'h10808, 'h108f7, 'h10818, 'h10828, 'h108f8, 'h10838, 'h10848, 'h108f9, 'h10af8, 'h103bc, 'h10858, 'h10868, 'h108fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h10878, 'h10888, 'h108fb, 'h10898, 'h108a8, 'h108fc, 'h108b8, 'h108c8, 'h108fd, 'h108d8, 'h106e8, 'h108fe, 'h10b08, 'h106f8, 'h103bc, 'h10708, 'h108ff, 'h10718, 'h21f8e, 'h21f8f, 'h21f8d, 'h10728, 'h10900, 'h10738, 'h10748, 'h10901, 'h10758, 'h10768, 'h10902, 'h10778, 'h10788, 'h10903, 'h10798, 'h10b08, 'h107a8, 'h10904, 'h103bc, 'h107b8, 'h107c8, 'h10905, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d8, 'h107e8, 'h10906, 'h107f8, 'h10808, 'h10907, 'h10818, 'h10828, 'h10908, 'h10838, 'h10848, 'h10909, 'h10b08, 'h10858, 'h103bc, 'h10868, 'h1090a, 'h10878, 'h21f8e, 'h21f8f, 'h21f8d, 'h10888, 'h1090b, 'h10898, 'h108a8, 'h1090c, 'h108b8, 'h108c8, 'h1090d, 'h108d8, 'h106e8, 'h1090e, 'h10b18, 'h106f8, 'h10708, 'h1090f, 'h103bc, 'h10718, 'h10728, 'h10910, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10748, 'h10911, 'h10758, 'h10768, 'h10912, 'h10778, 'h10788, 'h10913, 'h10798, 'h10b18, 'h107a8, 'h10914, 'h107b8, 'h103bc, 'h107c8, 'h10915, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e8, 'h10916, 'h107f8, 'h10808, 'h10917, 'h10818, 'h10828, 'h10918, 'h10838, 'h10848, 'h10919, 'h10b18, 'h10858, 'h10868, 'h1091a, 'h103bc, 'h10878, 'h10888, 'h1091b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10898, 'h108a8, 'h1091c, 'h108b8, 'h108c8, 'h1091d, 'h108d8, 'h106e8, 'h1091e, 'h10b28, 'h106f8, 'h10708, 'h1091f, 'h10718, 'h103bc, 'h10728, 'h10920, 'h10738, 'h21f8e, 'h21f8f, 'h21f8d, 'h10748, 'h10921, 'h10758, 'h10768, 'h10922, 'h10778, 'h10788, 'h10923, 'h10798, 'h10b28, 'h107a8, 'h10924, 'h107b8, 'h107c8, 'h10925, 'h103bc, 'h107d8, 'h107e8, 'h10926, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f8, 'h10808, 'h10927, 'h10818, 'h10828, 'h10928, 'h10838, 'h10848, 'h10929, 'h10b28, 'h10858, 'h10868, 'h1092a, 'h10878, 'h103bc, 'h10888, 'h1092b, 'h10898, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a8, 'h1092c, 'h108b8, 'h108c8, 'h1092d, 'h108d8, 'h106e8, 'h1092e, 'h10b38, 'h106f8, 'h10708, 'h1092f, 'h10718, 'h10728, 'h10930, 'h103bc, 'h10738, 'h10748, 'h10931, 'h21f8e, 'h21f8f, 'h21f8d, 'h10758, 'h10768, 'h10932, 'h10778, 'h10788, 'h10933, 'h10798, 'h10b38, 'h107a8, 'h10934, 'h107b8, 'h107c8, 'h10935, 'h107d8, 'h103bc, 'h107e8, 'h10936, 'h107f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10808, 'h10937, 'h10818, 'h10828, 'h10938, 'h10838, 'h10848, 'h10939, 'h10b38, 'h10858, 'h10868, 'h1093a, 'h10878, 'h10888, 'h1093b, 'h103bc, 'h10898, 'h108a8, 'h1093c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b8, 'h108c8, 'h1093d, 'h108d8, 'h106e8, 'h1093e, 'h10b48, 'h106f8, 'h10708, 'h1093f, 'h10718, 'h10728, 'h10940, 'h10738, 'h103bc, 'h10748, 'h10941, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h10768, 'h10942, 'h10778, 'h10788, 'h10943, 'h10798, 'h10b48, 'h107a8, 'h10944, 'h107b8, 'h107c8, 'h10945, 'h107d8, 'h107e8, 'h10946, 'h103bc, 'h107f8, 'h10808, 'h10947, 'h21f8e, 'h21f8f, 'h21f8d, 'h10818, 'h10828, 'h10948, 'h10838, 'h10848, 'h10949, 'h10b48, 'h10858, 'h10868, 'h1094a, 'h10878, 'h10888, 'h1094b, 'h10898, 'h103bc, 'h108a8, 'h1094c, 'h108b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c8, 'h1094d, 'h108d8, 'h106e8, 'h1094e, 'h10b58, 'h106f8, 'h10708, 'h1094f, 'h10718, 'h10728, 'h10950, 'h10738, 'h10748, 'h10951, 'h103bc, 'h10758, 'h10768, 'h10952, 'h21f8e, 'h21f8f, 'h21f8d, 'h10778, 'h10788, 'h10953, 'h10798, 'h10b58, 'h107a8, 'h10954, 'h107b8, 'h107c8, 'h10955, 'h107d8, 'h107e8, 'h10956, 'h107f8, 'h103bc, 'h10808, 'h10957, 'h10818, 'h21f8e, 'h21f8f, 'h21f8d, 'h10828, 'h10958, 'h10838, 'h10848, 'h10959, 'h10b58, 'h10858, 'h10868, 'h1095a, 'h10878, 'h10888, 'h1095b, 'h10898, 'h108a8, 'h1095c, 'h103bc, 'h108b8, 'h108c8, 'h1095d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d8, 'h106e8, 'h1095e, 'h10b68, 'h106f8, 'h10708, 'h1095f, 'h10718, 'h10728, 'h10960, 'h10738, 'h10748, 'h10961, 'h10758, 'h103bc, 'h10768, 'h10962, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10788, 'h10963, 'h10798, 'h10b68, 'h107a8, 'h10964, 'h107b8, 'h107c8, 'h10965, 'h107d8, 'h107e8, 'h10966, 'h107f8, 'h10808, 'h10967, 'h103bc, 'h10818, 'h10828, 'h10968, 'h21f8e, 'h21f8f, 'h21f8d, 'h10838, 'h10848, 'h10969, 'h10b68, 'h10858, 'h10868, 'h1096a, 'h10878, 'h10888, 'h1096b, 'h10898, 'h108a8, 'h1096c, 'h108b8, 'h103bc, 'h108c8, 'h1096d, 'h108d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e8, 'h1096e, 'h10b78, 'h106f8, 'h10708, 'h1096f, 'h10718, 'h10728, 'h10970, 'h10738, 'h10748, 'h10971, 'h10758, 'h10768, 'h10972, 'h103bc, 'h10778, 'h10788, 'h10973, 'h21f8e, 'h21f8f, 'h21f8d, 'h10798, 'h10b78, 'h107a8, 'h10974, 'h107b8, 'h107c8, 'h10975, 'h107d8, 'h107e8, 'h10976, 'h107f8, 'h10808, 'h10977, 'h10818, 'h103bc, 'h10828, 'h10978, 'h10838, 'h21f8e, 'h21f8f, 'h21f8d, 'h10848, 'h10979, 'h10b78, 'h10858, 'h10868, 'h1097a, 'h10878, 'h10888, 'h1097b, 'h10898, 'h108a8, 'h1097c, 'h108b8, 'h108c8, 'h1097d, 'h103bc, 'h108d8, 'h106e8, 'h1097e, 'h10b88, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f8, 'h10708, 'h1097f, 'h10718, 'h10728, 'h10980, 'h10738, 'h10748, 'h10981, 'h10758, 'h10768, 'h10982, 'h10778, 'h103bc, 'h10788, 'h10983, 'h10798, 'h10b88, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a8, 'h10984, 'h107b8, 'h107c8, 'h10985, 'h107d8, 'h107e8, 'h10986, 'h107f8, 'h10808, 'h10987, 'h10818, 'h10828, 'h10988, 'h103bc, 'h10838, 'h10848, 'h10989, 'h10b88, 'h21f8e, 'h21f8f, 'h21f8d, 'h10858, 'h10868, 'h1098a, 'h10878, 'h10888, 'h1098b, 'h10898, 'h108a8, 'h1098c, 'h108b8, 'h108c8, 'h1098d, 'h108d8, 'h103bc, 'h106e8, 'h1098e, 'h10b98, 'h106f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h1098f, 'h10718, 'h10728, 'h10990, 'h10738, 'h10748, 'h10991, 'h10758, 'h10768, 'h10992, 'h10778, 'h10788, 'h10993, 'h103bc, 'h10798, 'h10b98, 'h107a8, 'h10994, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b8, 'h107c8, 'h10995, 'h107d8, 'h107e8, 'h10996, 'h107f8, 'h10808, 'h10997, 'h10818, 'h10828, 'h10998, 'h10838, 'h103bc, 'h10848, 'h10999, 'h10b98, 'h10858, 'h21f8e, 'h21f8f, 'h21f8d, 'h10868, 'h1099a, 'h10878, 'h10888, 'h1099b, 'h10898, 'h108a8, 'h1099c, 'h108b8, 'h108c8, 'h1099d, 'h108d8, 'h106e8, 'h1099e, 'h10ba8, 'h103bc, 'h106f8, 'h10708, 'h1099f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10718, 'h10728, 'h109a0, 'h10738, 'h10748, 'h109a1, 'h10758, 'h10768, 'h109a2, 'h10778, 'h10788, 'h109a3, 'h10798, 'h10ba8, 'h103bc, 'h107a8, 'h109a4, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c8, 'h109a5, 'h107d8, 'h107e8, 'h109a6, 'h107f8, 'h10808, 'h109a7, 'h10818, 'h10828, 'h109a8, 'h10838, 'h10848, 'h109a9, 'h10ba8, 'h103bc, 'h10858, 'h10868, 'h109aa, 'h21f8e, 'h21f8f, 'h21f8d, 'h10878, 'h10888, 'h109ab, 'h10898, 'h108a8, 'h109ac, 'h108b8, 'h108c8, 'h109ad, 'h108d8, 'h106e8, 'h109ae, 'h10bb8, 'h106f8, 'h103bc, 'h10708, 'h109af, 'h10718, 'h21f8e, 'h21f8f, 'h21f8d, 'h10728, 'h109b0, 'h10738, 'h10748, 'h109b1, 'h10758, 'h10768, 'h109b2, 'h10778, 'h10788, 'h109b3, 'h10798, 'h10bb8, 'h107a8, 'h109b4, 'h103bc, 'h107b8, 'h107c8, 'h109b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d8, 'h107e8, 'h109b6, 'h107f8, 'h10808, 'h109b7, 'h10818, 'h10828, 'h109b8, 'h10838, 'h10848, 'h109b9, 'h10bb8, 'h10858, 'h103bc, 'h10868, 'h109ba, 'h10878, 'h21f8e, 'h21f8f, 'h21f8d, 'h10888, 'h109bb, 'h10898, 'h108a8, 'h109bc, 'h108b8, 'h108c8, 'h109bd, 'h108d8, 'h106e8, 'h109be, 'h10bc8, 'h106f8, 'h10708, 'h109bf, 'h103bc, 'h10718, 'h10728, 'h109c0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10748, 'h109c1, 'h10758, 'h10768, 'h109c2, 'h10778, 'h10788, 'h109c3, 'h10798, 'h10bc8, 'h107a8, 'h109c4, 'h107b8, 'h103bc, 'h107c8, 'h109c5, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e8, 'h109c6, 'h107f8, 'h10808, 'h109c7, 'h10818, 'h10828, 'h109c8, 'h10838, 'h10848, 'h109c9, 'h10bc8, 'h10858, 'h10868, 'h109ca, 'h103bc, 'h10878, 'h10888, 'h109cb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10898, 'h108a8, 'h109cc, 'h108b8, 'h108c8, 'h109cd, 'h108d8, 'h106e8, 'h109ce, 'h10bd8, 'h106f8, 'h10708, 'h109cf, 'h10718, 'h103bc, 'h10728, 'h109d0, 'h10738, 'h21f8e, 'h21f8f, 'h21f8d, 'h10748, 'h109d1, 'h10758, 'h10768, 'h109d2, 'h10778, 'h10788, 'h109d3, 'h10798, 'h10bd8, 'h107a8, 'h109d4, 'h107b8, 'h107c8, 'h109d5, 'h103bc, 'h107d8, 'h107e8, 'h109d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f8, 'h10808, 'h109d7, 'h10818, 'h10828, 'h109d8, 'h10838, 'h10848, 'h109d9, 'h10bd8, 'h10858, 'h10868, 'h109da, 'h10878, 'h103bc, 'h10888, 'h109db, 'h10898, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a8, 'h109dc, 'h108b8, 'h108c8, 'h109dd, 'h108d8, 'h106e8, 'h109de, 'h10be8, 'h106f8, 'h10708, 'h109df, 'h10718, 'h10728, 'h109e0, 'h103bc, 'h10738, 'h10748, 'h109e1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10758, 'h10768, 'h109e2, 'h10778, 'h10788, 'h109e3, 'h10798, 'h10be8, 'h107a8, 'h109e4, 'h107b8, 'h107c8, 'h109e5, 'h107d8, 'h103bc, 'h107e8, 'h109e6, 'h107f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10808, 'h109e7, 'h10818, 'h10828, 'h109e8, 'h10838, 'h10848, 'h109e9, 'h10be8, 'h10858, 'h10868, 'h109ea, 'h10878, 'h10888, 'h109eb, 'h103bc, 'h10898, 'h108a8, 'h109ec, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b8, 'h108c8, 'h109ed, 'h108d8, 'h106e8, 'h109ee, 'h10bf8, 'h106f8, 'h10708, 'h109ef, 'h10718, 'h10728, 'h109f0, 'h10738, 'h103bc, 'h10748, 'h109f1, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h10768, 'h109f2, 'h10778, 'h10788, 'h109f3, 'h10798, 'h10bf8, 'h107a8, 'h109f4, 'h107b8, 'h107c8, 'h109f5, 'h107d8, 'h107e8, 'h109f6, 'h103bc, 'h107f8, 'h10808, 'h109f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10818, 'h10828, 'h109f8, 'h10838, 'h10848, 'h109f9, 'h10bf8, 'h10858, 'h10868, 'h109fa, 'h10878, 'h10888, 'h109fb, 'h10898, 'h103bc, 'h108a8, 'h109fc, 'h108b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c8, 'h109fd, 'h108d8, 'h106e8, 'h109fe, 'h10c08, 'h106f8, 'h10708, 'h109ff, 'h10718, 'h10728, 'h10a00, 'h10738, 'h10748, 'h10a01, 'h103bc, 'h10758, 'h10768, 'h10a02, 'h21f8e, 'h21f8f, 'h21f8d, 'h10778, 'h10788, 'h10a03, 'h10798, 'h10c08, 'h107a8, 'h10a04, 'h107b8, 'h107c8, 'h10a05, 'h107d8, 'h107e8, 'h10a06, 'h107f8, 'h103bc, 'h10808, 'h10a07, 'h10818, 'h21f8e, 'h21f8f, 'h21f8d, 'h10828, 'h10a08, 'h10838, 'h10848, 'h10a09, 'h10c08, 'h10858, 'h10868, 'h10a0a, 'h10878, 'h10888, 'h10a0b, 'h10898, 'h108a8, 'h10a0c, 'h103bc, 'h108b8, 'h108c8, 'h10a0d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d8, 'h106e8, 'h10a0e, 'h10c18, 'h106f8, 'h10708, 'h10a0f, 'h10718, 'h10728, 'h10a10, 'h10738, 'h10748, 'h10a11, 'h10758, 'h103bc, 'h10768, 'h10a12, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10788, 'h10a13, 'h10798, 'h10c18, 'h107a8, 'h10a14, 'h107b8, 'h107c8, 'h10a15, 'h107d8, 'h107e8, 'h10a16, 'h107f8, 'h10808, 'h10a17, 'h103bc, 'h10818, 'h10828, 'h10a18, 'h21f8e, 'h21f8f, 'h21f8d, 'h10838, 'h10848, 'h10a19, 'h10c18, 'h10858, 'h10868, 'h10a1a, 'h10878, 'h10888, 'h10a1b, 'h10898, 'h108a8, 'h10a1c, 'h108b8, 'h103bc, 'h108c8, 'h10a1d, 'h108d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e8, 'h10a1e, 'h10c28, 'h106f8, 'h10708, 'h10a1f, 'h10718, 'h10728, 'h10a20, 'h10738, 'h10748, 'h10a21, 'h10758, 'h10768, 'h10a22, 'h103bc, 'h10778, 'h10788, 'h10a23, 'h21f8e, 'h21f8f, 'h21f8d, 'h10798, 'h10c28, 'h107a8, 'h10a24, 'h107b8, 'h107c8, 'h10a25, 'h107d8, 'h107e8, 'h10a26, 'h107f8, 'h10808, 'h10a27, 'h10818, 'h103bc, 'h10828, 'h10a28, 'h10838, 'h21f8e, 'h21f8f, 'h21f8d, 'h10848, 'h10a29, 'h10c28, 'h10858, 'h10868, 'h10a2a, 'h10878, 'h10888, 'h10a2b, 'h10898, 'h108a8, 'h10a2c, 'h108b8, 'h108c8, 'h10a2d, 'h103bc, 'h108d8, 'h106e8, 'h10a2e, 'h10c38, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f8, 'h10708, 'h10a2f, 'h10718, 'h10728, 'h10a30, 'h10738, 'h10748, 'h10a31, 'h10758, 'h10768, 'h10a32, 'h10778, 'h103bc, 'h10788, 'h10a33, 'h10798, 'h10c38, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a8, 'h10a34, 'h107b8, 'h107c8, 'h10a35, 'h107d8, 'h107e8, 'h10a36, 'h107f8, 'h10808, 'h10a37, 'h10818, 'h10828, 'h10a38, 'h103bc, 'h10838, 'h10848, 'h10a39, 'h10c38, 'h21f8e, 'h21f8f, 'h21f8d, 'h10858, 'h10868, 'h10a3a, 'h10878, 'h10888, 'h10a3b, 'h10898, 'h108a8, 'h10a3c, 'h108b8, 'h108c8, 'h10a3d, 'h108d8, 'h103bc, 'h106e8, 'h10a3e, 'h10c48, 'h106f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10a3f, 'h10718, 'h10728, 'h10a40, 'h10738, 'h10748, 'h10a41, 'h10758, 'h10768, 'h10a42, 'h10778, 'h10788, 'h10a43, 'h103bc, 'h10798, 'h10c48, 'h107a8, 'h10a44, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b8, 'h107c8, 'h10a45, 'h107d8, 'h107e8, 'h10a46, 'h107f8, 'h10808, 'h10a47, 'h10818, 'h10828, 'h10a48, 'h10838, 'h103bc, 'h10848, 'h10a49, 'h10c48, 'h10858, 'h21f8e, 'h21f8f, 'h21f8d, 'h10868, 'h10a4a, 'h10878, 'h10888, 'h10a4b, 'h10898, 'h108a8, 'h10a4c, 'h108b8, 'h108c8, 'h10a4d, 'h108d8, 'h106e8, 'h10a4e, 'h10c58, 'h103bc, 'h106f8, 'h10708, 'h10a4f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10718, 'h10728, 'h10a50, 'h10738, 'h10748, 'h10a51, 'h10758, 'h10768, 'h10a52, 'h10778, 'h10788, 'h10a53, 'h10798, 'h10c58, 'h103bc, 'h107a8, 'h10a54, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c8, 'h10a55, 'h107d8, 'h107e8, 'h10a56, 'h107f8, 'h10808, 'h10a57, 'h10818, 'h10828, 'h10a58, 'h10838, 'h10848, 'h10a59, 'h10c58, 'h103bc, 'h10858, 'h10868, 'h10a5a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10878, 'h10888, 'h10a5b, 'h10898, 'h108a8, 'h10a5c, 'h108b8, 'h108c8, 'h10a5d, 'h108d8, 'h106e8, 'h10a5e, 'h10c68, 'h106f8, 'h103bc, 'h10708, 'h10a5f, 'h10718, 'h21f8e, 'h21f8f, 'h21f8d, 'h10728, 'h10a60, 'h10738, 'h10748, 'h10a61, 'h10758, 'h10768, 'h10a62, 'h10778, 'h10788, 'h10a63, 'h10798, 'h10c68, 'h107a8, 'h10a64, 'h103bc, 'h107b8, 'h107c8, 'h10a65, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d8, 'h107e8, 'h10a66, 'h107f8, 'h10808, 'h10a67, 'h10818, 'h10828, 'h10a68, 'h10838, 'h10848, 'h10a69, 'h10c68, 'h10858, 'h103bc, 'h10868, 'h10a6a, 'h10878, 'h21f8e, 'h21f8f, 'h21f8d, 'h10888, 'h10a6b, 'h10898, 'h108a8, 'h10a6c, 'h108b8, 'h108c8, 'h10a6d, 'h108d8, 'h106e8, 'h10a6e, 'h10c78, 'h106f8, 'h10708, 'h10a6f, 'h103bc, 'h10718, 'h10728, 'h10a70, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10748, 'h10a71, 'h10758, 'h10768, 'h10a72, 'h10778, 'h10788, 'h10a73, 'h10798, 'h10c78, 'h107a8, 'h10a74, 'h107b8, 'h103bc, 'h107c8, 'h10a75, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e8, 'h10a76, 'h107f8, 'h10808, 'h10a77, 'h10818, 'h10828, 'h10a78, 'h10838, 'h10848, 'h10a79, 'h10c78, 'h10858, 'h10868, 'h10a7a, 'h103bc, 'h10878, 'h10888, 'h10a7b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10898, 'h108a8, 'h10a7c, 'h108b8, 'h108c8, 'h10a7d, 'h108d8, 'h106e8, 'h10a7e, 'h10c88, 'h106f8, 'h10708, 'h10a7f, 'h10718, 'h103bc, 'h10728, 'h10a80, 'h10738, 'h21f8e, 'h21f8f, 'h21f8d, 'h10748, 'h10a81, 'h10758, 'h10768, 'h10a82, 'h10778, 'h10788, 'h10a83, 'h10798, 'h10c88, 'h107a8, 'h10a84, 'h107b8, 'h107c8, 'h10a85, 'h103bc, 'h107d8, 'h107e8, 'h10a86, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f8, 'h10808, 'h10a87, 'h10818, 'h10828, 'h10a88, 'h10838, 'h10848, 'h10a89, 'h10c88, 'h10858, 'h10868, 'h10a8a, 'h10878, 'h103bc, 'h10888, 'h10a8b, 'h10898, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a8, 'h10a8c, 'h108b8, 'h108c8, 'h10a8d, 'h108d8, 'h106e8, 'h10a8e, 'h10c98, 'h106f8, 'h10708, 'h10a8f, 'h10718, 'h10728, 'h10a90, 'h103bc, 'h10738, 'h10748, 'h10a91, 'h21f8e, 'h21f8f, 'h21f8d, 'h10758, 'h10768, 'h10a92, 'h10778, 'h10788, 'h10a93, 'h10798, 'h10c98, 'h107a8, 'h10a94, 'h107b8, 'h107c8, 'h10a95, 'h107d8, 'h103bc, 'h107e8, 'h10a96, 'h107f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10808, 'h10a97, 'h10818, 'h10828, 'h10a98, 'h10838, 'h10848, 'h10a99, 'h10c98, 'h10858, 'h10868, 'h10a9a, 'h10878, 'h10888, 'h10a9b, 'h103bc, 'h10898, 'h108a8, 'h10a9c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b8, 'h108c8, 'h10a9d, 'h108d8, 'h106e8, 'h10a9e, 'h10ca8, 'h106f8, 'h10708, 'h10a9f, 'h10718, 'h10728, 'h10aa0, 'h10738, 'h103bc, 'h10748, 'h10aa1, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h10768, 'h10aa2, 'h10778, 'h10788, 'h10aa3, 'h10798, 'h10ca8, 'h107a8, 'h10aa4, 'h107b8, 'h107c8, 'h10aa5, 'h107d8, 'h107e8, 'h10aa6, 'h103bc, 'h107f8, 'h10808, 'h10aa7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10818, 'h10828, 'h10aa8, 'h10838, 'h10848, 'h10aa9, 'h10ca8, 'h10858, 'h10868, 'h10aaa, 'h10878, 'h10888, 'h10aab, 'h10898, 'h103bc, 'h108a8, 'h10aac, 'h108b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c8, 'h10aad, 'h108d8, 'h106e8, 'h10aae, 'h10cb8, 'h106f8, 'h10708, 'h10aaf, 'h10718, 'h10728, 'h10ab0, 'h10738, 'h10748, 'h10ab1, 'h103bc, 'h10758, 'h10768, 'h10ab2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10778, 'h10788, 'h10ab3, 'h10798, 'h10cb8, 'h107a8, 'h10ab4, 'h107b8, 'h107c8, 'h10ab5, 'h107d8, 'h107e8, 'h10ab6, 'h107f8, 'h103bc, 'h10808, 'h10ab7, 'h10818, 'h21f8e, 'h21f8f, 'h21f8d, 'h10828, 'h10ab8, 'h10838, 'h10848, 'h10ab9, 'h10cb8, 'h10858, 'h10868, 'h10aba, 'h10878, 'h10888, 'h10abb, 'h10898, 'h108a8, 'h10abc, 'h103bc, 'h108b8, 'h108c8, 'h10abd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d8, 'h106e8, 'h10abe, 'h10cc8, 'h106f8, 'h10708, 'h10abf, 'h10718, 'h10728, 'h10ac0, 'h10738, 'h10748, 'h10ac1, 'h10758, 'h103bc, 'h10768, 'h10ac2, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10788, 'h10ac3, 'h10798, 'h10cc8, 'h107a8, 'h10ac4, 'h107b8, 'h107c8, 'h10ac5, 'h107d8, 'h107e8, 'h10ac6, 'h107f8, 'h10808, 'h10ac7, 'h103bc, 'h10818, 'h10828, 'h10ac8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10838, 'h10848, 'h10ac9, 'h10cc8, 'h10858, 'h10868, 'h10aca, 'h10878, 'h10888, 'h10acb, 'h10898, 'h108a8, 'h10acc, 'h108b8, 'h103bc, 'h108c8, 'h10acd, 'h108d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e8, 'h10ace, 'h10cd8, 'h106f8, 'h10708, 'h10acf, 'h10718, 'h10728, 'h10ad0, 'h10738, 'h10748, 'h10ad1, 'h10758, 'h10768, 'h10ad2, 'h103bc, 'h10778, 'h10788, 'h10ad3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10798, 'h10cd8, 'h107a8, 'h10ad4, 'h107b8, 'h107c8, 'h10ad5, 'h107d8, 'h107e8, 'h10ad6, 'h107f8, 'h10808, 'h10ad7, 'h10818, 'h103bc, 'h10828, 'h10ad8, 'h10838, 'h21f8e, 'h21f8f, 'h21f8d, 'h10848, 'h10ad9, 'h10cd8, 'h10858, 'h10868, 'h10ada, 'h10878, 'h10888, 'h10adb, 'h10898, 'h108a8, 'h10adc, 'h108b8, 'h108c8, 'h10add, 'h103bc, 'h108d8, 'h106e8, 'h108de, 'h10ae8, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f8, 'h10708, 'h108df, 'h10718, 'h10728, 'h108e0, 'h10738, 'h10748, 'h108e1, 'h10758, 'h10768, 'h108e2, 'h10778, 'h103bc, 'h10788, 'h108e3, 'h10798, 'h10ae8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a8, 'h108e4, 'h107b8, 'h107c8, 'h108e5, 'h107d8, 'h107e8, 'h108e6, 'h107f8, 'h10808, 'h108e7, 'h10818, 'h10828, 'h108e8, 'h103bc, 'h10838, 'h10848, 'h108e9, 'h10ae8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10858, 'h10868, 'h108ea, 'h10878, 'h10888, 'h108eb, 'h10898, 'h108a8, 'h108ec, 'h108b8, 'h108c8, 'h108ed, 'h108d8, 'h103bc, 'h106e8, 'h108ee, 'h10af8, 'h106f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h108ef, 'h10718, 'h10728, 'h108f0, 'h10738, 'h10748, 'h108f1, 'h10758, 'h10768, 'h108f2, 'h10778, 'h10788, 'h108f3, 'h103bc, 'h10798, 'h10af8, 'h107a8, 'h108f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b8, 'h107c8, 'h108f5, 'h107d8, 'h107e8, 'h108f6, 'h107f8, 'h10808, 'h108f7, 'h10818, 'h10828, 'h108f8, 'h10838, 'h103bc, 'h10848, 'h108f9, 'h10af8, 'h10858, 'h21f8e, 'h21f8f, 'h21f8d, 'h10868, 'h108fa, 'h10878, 'h10888, 'h108fb, 'h10898, 'h108a8, 'h108fc, 'h108b8, 'h108c8, 'h108fd, 'h108d8, 'h106e8, 'h108fe, 'h10b08, 'h103bc, 'h106f8, 'h10708, 'h108ff, 'h21f8e, 'h21f8f, 'h21f8d, 'h10718, 'h10728, 'h10900, 'h10738, 'h10748, 'h10901, 'h10758, 'h10768, 'h10902, 'h10778, 'h10788, 'h10903, 'h10798, 'h10b08, 'h103bc, 'h107a8, 'h10904, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c8, 'h10905, 'h107d8, 'h107e8, 'h10906, 'h107f8, 'h10808, 'h10907, 'h10818, 'h10828, 'h10908, 'h10838, 'h10848, 'h10909, 'h10b08, 'h103bc, 'h10858, 'h10868, 'h1090a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10878, 'h10888, 'h1090b, 'h10898, 'h108a8, 'h1090c, 'h108b8, 'h108c8, 'h1090d, 'h108d8, 'h106e8, 'h1090e, 'h10b18, 'h106f8, 'h103bc, 'h10708, 'h1090f, 'h10718, 'h21f8e, 'h21f8f, 'h21f8d, 'h10728, 'h10910, 'h10738, 'h10748, 'h10911, 'h10758, 'h10768, 'h10912, 'h10778, 'h10788, 'h10913, 'h10798, 'h10b18, 'h107a8, 'h10914, 'h103bc, 'h107b8, 'h107c8, 'h10915, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d8, 'h107e8, 'h10916, 'h107f8, 'h10808, 'h10917, 'h10818, 'h10828, 'h10918, 'h10838, 'h10848, 'h10919, 'h10b18, 'h10858, 'h103bc, 'h10868, 'h1091a, 'h10878, 'h21f8e, 'h21f8f, 'h21f8d, 'h10888, 'h1091b, 'h10898, 'h108a8, 'h1091c, 'h108b8, 'h108c8, 'h1091d, 'h108d8, 'h106e8, 'h1091e, 'h10b28, 'h106f8, 'h10708, 'h1091f, 'h103bc, 'h10718, 'h10728, 'h10920, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10748, 'h10921, 'h10758, 'h10768, 'h10922, 'h10778, 'h10788, 'h10923, 'h10798, 'h10b28, 'h107a8, 'h10924, 'h107b8, 'h103bc, 'h107c8, 'h10925, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e8, 'h10926, 'h107f8, 'h10808, 'h10927, 'h10818, 'h10828, 'h10928, 'h10838, 'h10848, 'h10929, 'h10b28, 'h10858, 'h10868, 'h1092a, 'h103bc, 'h10878, 'h10888, 'h1092b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10898, 'h108a8, 'h1092c, 'h108b8, 'h108c8, 'h1092d, 'h108d8, 'h106e8, 'h1092e, 'h10b38, 'h106f8, 'h10708, 'h1092f, 'h10718, 'h103bc, 'h10728, 'h10930, 'h10738, 'h21f8e, 'h21f8f, 'h21f8d, 'h10748, 'h10931, 'h10758, 'h10768, 'h10932, 'h10778, 'h10788, 'h10933, 'h10798, 'h10b38, 'h107a8, 'h10934, 'h107b8, 'h107c8, 'h10935, 'h103bc, 'h107d8, 'h107e8, 'h10936, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f8, 'h10808, 'h10937, 'h10818, 'h10828, 'h10938, 'h10838, 'h10848, 'h10939, 'h10b38, 'h10858, 'h10868, 'h1093a, 'h10878, 'h103bc, 'h10888, 'h1093b, 'h10898, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a8, 'h1093c, 'h108b8, 'h108c8, 'h1093d, 'h108d8, 'h106e8, 'h1093e, 'h10b48, 'h106f8, 'h10708, 'h1093f, 'h10718, 'h10728, 'h10940, 'h103bc, 'h10738, 'h10748, 'h10941, 'h21f8e, 'h21f8f, 'h21f8d, 'h10758, 'h10768, 'h10942, 'h10778, 'h10788, 'h10943, 'h10798, 'h10b48, 'h107a8, 'h10944, 'h107b8, 'h107c8, 'h10945, 'h107d8, 'h103bc, 'h107e8, 'h10946, 'h107f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10808, 'h10947, 'h10818, 'h10828, 'h10948, 'h10838, 'h10848, 'h10949, 'h10b48, 'h10858, 'h10868, 'h1094a, 'h10878, 'h10888, 'h1094b, 'h103bc, 'h10898, 'h108a8, 'h1094c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b8, 'h108c8, 'h1094d, 'h108d8, 'h106e8, 'h1094e, 'h10b58, 'h106f8, 'h10708, 'h1094f, 'h10718, 'h10728, 'h10950, 'h10738, 'h103bc, 'h10748, 'h10951, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h10768, 'h10952, 'h10778, 'h10788, 'h10953, 'h10798, 'h10b58, 'h107a8, 'h10954, 'h107b8, 'h107c8, 'h10955, 'h107d8, 'h107e8, 'h10956, 'h103bc, 'h107f8, 'h10808, 'h10957, 'h21f8e, 'h21f8f, 'h21f8d, 'h10818, 'h10828, 'h10958, 'h10838, 'h10848, 'h10959, 'h10b58, 'h10858, 'h10868, 'h1095a, 'h10878, 'h10888, 'h1095b, 'h10898, 'h103bc, 'h108a8, 'h1095c, 'h108b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c8, 'h1095d, 'h108d8, 'h106e8, 'h1095e, 'h10b68, 'h106f8, 'h10708, 'h1095f, 'h10718, 'h10728, 'h10960, 'h10738, 'h10748, 'h10961, 'h103bc, 'h10758, 'h10768, 'h10962, 'h21f8e, 'h21f8f, 'h21f8d, 'h10778, 'h10788, 'h10963, 'h10798, 'h10b68, 'h107a8, 'h10964, 'h107b8, 'h107c8, 'h10965, 'h107d8, 'h107e8, 'h10966, 'h107f8, 'h103bc, 'h10808, 'h10967, 'h10818, 'h21f8e, 'h21f8f, 'h21f8d, 'h10828, 'h10968, 'h10838, 'h10848, 'h10969, 'h10b68, 'h10858, 'h10868, 'h1096a, 'h10878, 'h10888, 'h1096b, 'h10898, 'h108a8, 'h1096c, 'h103bc, 'h108b8, 'h108c8, 'h1096d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d8, 'h106e8, 'h1096e, 'h10b78, 'h106f8, 'h10708, 'h1096f, 'h10718, 'h10728, 'h10970, 'h10738, 'h10748, 'h10971, 'h10758, 'h103bc, 'h10768, 'h10972, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10788, 'h10973, 'h10798, 'h10b78, 'h107a8, 'h10974, 'h107b8, 'h107c8, 'h10975, 'h107d8, 'h107e8, 'h10976, 'h107f8, 'h10808, 'h10977, 'h103bc, 'h10818, 'h10828, 'h10978, 'h21f8e, 'h21f8f, 'h21f8d, 'h10838, 'h10848, 'h10979, 'h10b78, 'h10858, 'h10868, 'h1097a, 'h10878, 'h10888, 'h1097b, 'h10898, 'h108a8, 'h1097c, 'h108b8, 'h103bc, 'h108c8, 'h1097d, 'h108d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e8, 'h1097e, 'h10b88, 'h106f8, 'h10708, 'h1097f, 'h10718, 'h10728, 'h10980, 'h10738, 'h10748, 'h10981, 'h10758, 'h10768, 'h10982, 'h103bc, 'h10778, 'h10788, 'h10983, 'h21f8e, 'h21f8f, 'h21f8d, 'h10798, 'h10b88, 'h107a8, 'h10984, 'h107b8, 'h107c8, 'h10985, 'h107d8, 'h107e8, 'h10986, 'h107f8, 'h10808, 'h10987, 'h10818, 'h103bc, 'h10828, 'h10988, 'h10838, 'h21f8e, 'h21f8f, 'h21f8d, 'h10848, 'h10989, 'h10b88, 'h10858, 'h10868, 'h1098a, 'h10878, 'h10888, 'h1098b, 'h10898, 'h108a8, 'h1098c, 'h108b8, 'h108c8, 'h1098d, 'h103bc, 'h108d8, 'h106e8, 'h1098e, 'h10b98, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f8, 'h10708, 'h1098f, 'h10718, 'h10728, 'h10990, 'h10738, 'h10748, 'h10991, 'h10758, 'h10768, 'h10992, 'h10778, 'h103bc, 'h10788, 'h10993, 'h10798, 'h10b98, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a8, 'h10994, 'h107b8, 'h107c8, 'h10995, 'h107d8, 'h107e8, 'h10996, 'h107f8, 'h10808, 'h10997, 'h10818, 'h10828, 'h10998, 'h103bc, 'h10838, 'h10848, 'h10999, 'h10b98, 'h21f8e, 'h21f8f, 'h21f8d, 'h10858, 'h10868, 'h1099a, 'h10878, 'h10888, 'h1099b, 'h10898, 'h108a8, 'h1099c, 'h108b8, 'h108c8, 'h1099d, 'h108d8, 'h103bc, 'h106e8, 'h1099e, 'h10ba8, 'h106f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h1099f, 'h10718, 'h10728, 'h109a0, 'h10738, 'h10748, 'h109a1, 'h10758, 'h10768, 'h109a2, 'h10778, 'h10788, 'h109a3, 'h103bc, 'h10798, 'h10ba8, 'h107a8, 'h109a4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b8, 'h107c8, 'h109a5, 'h107d8, 'h107e8, 'h109a6, 'h107f8, 'h10808, 'h109a7, 'h10818, 'h10828, 'h109a8, 'h10838, 'h103bc, 'h10848, 'h109a9, 'h10ba8, 'h10858, 'h21f8e, 'h21f8f, 'h21f8d, 'h10868, 'h109aa, 'h10878, 'h10888, 'h109ab, 'h10898, 'h108a8, 'h109ac, 'h108b8, 'h108c8, 'h109ad, 'h108d8, 'h106e8, 'h109ae, 'h10bb8, 'h103bc, 'h106f8, 'h10708, 'h109af, 'h21f8e, 'h21f8f, 'h21f8d, 'h10718, 'h10728, 'h109b0, 'h10738, 'h10748, 'h109b1, 'h10758, 'h10768, 'h109b2, 'h10778, 'h10788, 'h109b3, 'h10798, 'h10bb8, 'h103bc, 'h107a8, 'h109b4, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c8, 'h109b5, 'h107d8, 'h107e8, 'h109b6, 'h107f8, 'h10808, 'h109b7, 'h10818, 'h10828, 'h109b8, 'h10838, 'h10848, 'h109b9, 'h10bb8, 'h103bc, 'h10858, 'h10868, 'h109ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h10878, 'h10888, 'h109bb, 'h10898, 'h108a8, 'h109bc, 'h108b8, 'h108c8, 'h109bd, 'h108d8, 'h106e8, 'h109be, 'h10bc8, 'h106f8, 'h103bc, 'h10708, 'h109bf, 'h10718, 'h21f8e, 'h21f8f, 'h21f8d, 'h10728, 'h109c0, 'h10738, 'h10748, 'h109c1, 'h10758, 'h10768, 'h109c2, 'h10778, 'h10788, 'h109c3, 'h10798, 'h10bc8, 'h107a8, 'h109c4, 'h103bc, 'h107b8, 'h107c8, 'h109c5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d8, 'h107e8, 'h109c6, 'h107f8, 'h10808, 'h109c7, 'h10818, 'h10828, 'h109c8, 'h10838, 'h10848, 'h109c9, 'h10bc8, 'h10858, 'h103bc, 'h10868, 'h109ca, 'h10878, 'h21f8e, 'h21f8f, 'h21f8d, 'h10888, 'h109cb, 'h10898, 'h108a8, 'h109cc, 'h108b8, 'h108c8, 'h109cd, 'h108d8, 'h106e8, 'h109ce, 'h10bd8, 'h106f8, 'h10708, 'h109cf, 'h103bc, 'h10718, 'h10728, 'h109d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10748, 'h109d1, 'h10758, 'h10768, 'h109d2, 'h10778, 'h10788, 'h109d3, 'h10798, 'h10bd8, 'h107a8, 'h109d4, 'h107b8, 'h103bc, 'h107c8, 'h109d5, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e8, 'h109d6, 'h107f8, 'h10808, 'h109d7, 'h10818, 'h10828, 'h109d8, 'h10838, 'h10848, 'h109d9, 'h10bd8, 'h10858, 'h10868, 'h109da, 'h103bc, 'h10878, 'h10888, 'h109db, 'h21f8e, 'h21f8f, 'h21f8d, 'h10898, 'h108a8, 'h109dc, 'h108b8, 'h108c8, 'h109dd, 'h108d8, 'h106e8, 'h109de, 'h10be8, 'h106f8, 'h10708, 'h109df, 'h10718, 'h103bc, 'h10728, 'h109e0, 'h10738, 'h21f8e, 'h21f8f, 'h21f8d, 'h10748, 'h109e1, 'h10758, 'h10768, 'h109e2, 'h10778, 'h10788, 'h109e3, 'h10798, 'h10be8, 'h107a8, 'h109e4, 'h107b8, 'h107c8, 'h109e5, 'h103bc, 'h107d8, 'h107e8, 'h109e6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f8, 'h10808, 'h109e7, 'h10818, 'h10828, 'h109e8, 'h10838, 'h10848, 'h109e9, 'h10be8, 'h10858, 'h10868, 'h109ea, 'h10878, 'h103bc, 'h10888, 'h109eb, 'h10898, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a8, 'h109ec, 'h108b8, 'h108c8, 'h109ed, 'h108d8, 'h106e8, 'h109ee, 'h10bf8, 'h106f8, 'h10708, 'h109ef, 'h10718, 'h10728, 'h109f0, 'h103bc, 'h10738, 'h10748, 'h109f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10758, 'h10768, 'h109f2, 'h10778, 'h10788, 'h109f3, 'h10798, 'h10bf8, 'h107a8, 'h109f4, 'h107b8, 'h107c8, 'h109f5, 'h107d8, 'h103bc, 'h107e8, 'h109f6, 'h107f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10808, 'h109f7, 'h10818, 'h10828, 'h109f8, 'h10838, 'h10848, 'h109f9, 'h10bf8, 'h10858, 'h10868, 'h109fa, 'h10878, 'h10888, 'h109fb, 'h103bc, 'h10898, 'h108a8, 'h109fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b8, 'h108c8, 'h109fd, 'h108d8, 'h106e8, 'h109fe, 'h10c08, 'h106f8, 'h10708, 'h109ff, 'h10718, 'h10728, 'h10a00, 'h10738, 'h103bc, 'h10748, 'h10a01, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h10768, 'h10a02, 'h10778, 'h10788, 'h10a03, 'h10798, 'h10c08, 'h107a8, 'h10a04, 'h107b8, 'h107c8, 'h10a05, 'h107d8, 'h107e8, 'h10a06, 'h103bc, 'h107f8, 'h10808, 'h10a07, 'h21f8e, 'h21f8f, 'h21f8d, 'h10818, 'h10828, 'h10a08, 'h10838, 'h10848, 'h10a09, 'h10c08, 'h10858, 'h10868, 'h10a0a, 'h10878, 'h10888, 'h10a0b, 'h10898, 'h103bc, 'h108a8, 'h10a0c, 'h108b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c8, 'h10a0d, 'h108d8, 'h106e8, 'h10a0e, 'h10c18, 'h106f8, 'h10708, 'h10a0f, 'h10718, 'h10728, 'h10a10, 'h10738, 'h10748, 'h10a11, 'h103bc, 'h10758, 'h10768, 'h10a12, 'h21f8e, 'h21f8f, 'h21f8d, 'h10778, 'h10788, 'h10a13, 'h10798, 'h10c18, 'h107a8, 'h10a14, 'h107b8, 'h107c8, 'h10a15, 'h107d8, 'h107e8, 'h10a16, 'h107f8, 'h103bc, 'h10808, 'h10a17, 'h10818, 'h21f8e, 'h21f8f, 'h21f8d, 'h10828, 'h10a18, 'h10838, 'h10848, 'h10a19, 'h10c18, 'h10858, 'h10868, 'h10a1a, 'h10878, 'h10888, 'h10a1b, 'h10898, 'h108a8, 'h10a1c, 'h103bc, 'h108b8, 'h108c8, 'h10a1d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d8, 'h106e8, 'h10a1e, 'h10c28, 'h106f8, 'h10708, 'h10a1f, 'h10718, 'h10728, 'h10a20, 'h10738, 'h10748, 'h10a21, 'h10758, 'h103bc, 'h10768, 'h10a22, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10788, 'h10a23, 'h10798, 'h10c28, 'h107a8, 'h10a24, 'h107b8, 'h107c8, 'h10a25, 'h107d8, 'h107e8, 'h10a26, 'h107f8, 'h10808, 'h10a27, 'h103bc, 'h10818, 'h10828, 'h10a28, 'h21f8e, 'h21f8f, 'h21f8d, 'h10838, 'h10848, 'h10a29, 'h10c28, 'h10858, 'h10868, 'h10a2a, 'h10878, 'h10888, 'h10a2b, 'h10898, 'h108a8, 'h10a2c, 'h108b8, 'h103bc, 'h108c8, 'h10a2d, 'h108d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e8, 'h10a2e, 'h10c38, 'h106f8, 'h10708, 'h10a2f, 'h10718, 'h10728, 'h10a30, 'h10738, 'h10748, 'h10a31, 'h10758, 'h10768, 'h10a32, 'h103bc, 'h10778, 'h10788, 'h10a33, 'h21f8e, 'h21f8f, 'h21f8d, 'h10798, 'h10c38, 'h107a8, 'h10a34, 'h107b8, 'h107c8, 'h10a35, 'h107d8, 'h107e8, 'h10a36, 'h107f8, 'h10808, 'h10a37, 'h10818, 'h103bc, 'h10828, 'h10a38, 'h10838, 'h21f8e, 'h21f8f, 'h21f8d, 'h10848, 'h10a39, 'h10c38, 'h10858, 'h10868, 'h10a3a, 'h10878, 'h10888, 'h10a3b, 'h10898, 'h108a8, 'h10a3c, 'h108b8, 'h108c8, 'h10a3d, 'h103bc, 'h108d8, 'h106e8, 'h10a3e, 'h10c48, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f8, 'h10708, 'h10a3f, 'h10718, 'h10728, 'h10a40, 'h10738, 'h10748, 'h10a41, 'h10758, 'h10768, 'h10a42, 'h10778, 'h103bc, 'h10788, 'h10a43, 'h10798, 'h10c48, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a8, 'h10a44, 'h107b8, 'h107c8, 'h10a45, 'h107d8, 'h107e8, 'h10a46, 'h107f8, 'h10808, 'h10a47, 'h10818, 'h10828, 'h10a48, 'h103bc, 'h10838, 'h10848, 'h10a49, 'h10c48, 'h21f8e, 'h21f8f, 'h21f8d, 'h10858, 'h10868, 'h10a4a, 'h10878, 'h10888, 'h10a4b, 'h10898, 'h108a8, 'h10a4c, 'h108b8, 'h108c8, 'h10a4d, 'h108d8, 'h103bc, 'h106e8, 'h10a4e, 'h10c58, 'h106f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10a4f, 'h10718, 'h10728, 'h10a50, 'h10738, 'h10748, 'h10a51, 'h10758, 'h10768, 'h10a52, 'h10778, 'h10788, 'h10a53, 'h103bc, 'h10798, 'h10c58, 'h107a8, 'h10a54, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b8, 'h107c8, 'h10a55, 'h107d8, 'h107e8, 'h10a56, 'h107f8, 'h10808, 'h10a57, 'h10818, 'h10828, 'h10a58, 'h10838, 'h103bc, 'h10848, 'h10a59, 'h10c58, 'h10858, 'h21f8e, 'h21f8f, 'h21f8d, 'h10868, 'h10a5a, 'h10878, 'h10888, 'h10a5b, 'h10898, 'h108a8, 'h10a5c, 'h108b8, 'h108c8, 'h10a5d, 'h108d8, 'h106e8, 'h10a5e, 'h10c68, 'h103bc, 'h106f8, 'h10708, 'h10a5f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10718, 'h10728, 'h10a60, 'h10738, 'h10748, 'h10a61, 'h10758, 'h10768, 'h10a62, 'h10778, 'h10788, 'h10a63, 'h10798, 'h10c68, 'h103bc, 'h107a8, 'h10a64, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c8, 'h10a65, 'h107d8, 'h107e8, 'h10a66, 'h107f8, 'h10808, 'h10a67, 'h10818, 'h10828, 'h10a68, 'h10838, 'h10848, 'h10a69, 'h10c68, 'h103bc, 'h10858, 'h10868, 'h10a6a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10878, 'h10888, 'h10a6b, 'h10898, 'h108a8, 'h10a6c, 'h108b8, 'h108c8, 'h10a6d, 'h108d8, 'h106e8, 'h10a6e, 'h10c78, 'h106f8, 'h103bc, 'h10708, 'h10a6f, 'h10718, 'h21f8e, 'h21f8f, 'h21f8d, 'h10728, 'h10a70, 'h10738, 'h10748, 'h10a71, 'h10758, 'h10768, 'h10a72, 'h10778, 'h10788, 'h10a73, 'h10798, 'h10c78, 'h107a8, 'h10a74, 'h103bc, 'h107b8, 'h107c8, 'h10a75, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d8, 'h107e8, 'h10a76, 'h107f8, 'h10808, 'h10a77, 'h10818, 'h10828, 'h10a78, 'h10838, 'h10848, 'h10a79, 'h10c78, 'h10858, 'h103bc, 'h10868, 'h10a7a, 'h10878, 'h21f8e, 'h21f8f, 'h21f8d, 'h10888, 'h10a7b, 'h10898, 'h108a8, 'h10a7c, 'h108b8, 'h108c8, 'h10a7d, 'h108d8, 'h106e8, 'h10a7e, 'h10c88, 'h106f8, 'h10708, 'h10a7f, 'h103bc, 'h10718, 'h10728, 'h10a80, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10748, 'h10a81, 'h10758, 'h10768, 'h10a82, 'h10778, 'h10788, 'h10a83, 'h10798, 'h10c88, 'h107a8, 'h10a84, 'h107b8, 'h103bc, 'h107c8, 'h10a85, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e8, 'h10a86, 'h107f8, 'h10808, 'h10a87, 'h10818, 'h10828, 'h10a88, 'h10838, 'h10848, 'h10a89, 'h10c88, 'h10858, 'h10868, 'h10a8a, 'h103bc, 'h10878, 'h10888, 'h10a8b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10898, 'h108a8, 'h10a8c, 'h108b8, 'h108c8, 'h10a8d, 'h108d8, 'h106e8, 'h10a8e, 'h10c98, 'h106f8, 'h10708, 'h10a8f, 'h10718, 'h103bc, 'h10728, 'h10a90, 'h10738, 'h21f8e, 'h21f8f, 'h21f8d, 'h10748, 'h10a91, 'h10758, 'h10768, 'h10a92, 'h10778, 'h10788, 'h10a93, 'h10798, 'h10c98, 'h107a8, 'h10a94, 'h107b8, 'h107c8, 'h10a95, 'h103bc, 'h107d8, 'h107e8, 'h10a96, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f8, 'h10808, 'h10a97, 'h10818, 'h10828, 'h10a98, 'h10838, 'h10848, 'h10a99, 'h10c98, 'h10858, 'h10868, 'h10a9a, 'h10878, 'h103bc, 'h10888, 'h10a9b, 'h10898, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a8, 'h10a9c, 'h108b8, 'h108c8, 'h10a9d, 'h108d8, 'h106e8, 'h10a9e, 'h10ca8, 'h106f8, 'h10708, 'h10a9f, 'h10718, 'h10728, 'h10aa0, 'h103bc, 'h10738, 'h10748, 'h10aa1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10758, 'h10768, 'h10aa2, 'h10778, 'h10788, 'h10aa3, 'h10798, 'h10ca8, 'h107a8, 'h10aa4, 'h107b8, 'h107c8, 'h10aa5, 'h107d8, 'h103bc, 'h107e8, 'h10aa6, 'h107f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10808, 'h10aa7, 'h10818, 'h10828, 'h10aa8, 'h10838, 'h10848, 'h10aa9, 'h10ca8, 'h10858, 'h10868, 'h10aaa, 'h10878, 'h10888, 'h10aab, 'h103bc, 'h10898, 'h108a8, 'h10aac, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b8, 'h108c8, 'h10aad, 'h108d8, 'h106e8, 'h10aae, 'h10cb8, 'h106f8, 'h10708, 'h10aaf, 'h10718, 'h10728, 'h10ab0, 'h10738, 'h103bc, 'h10748, 'h10ab1, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h10768, 'h10ab2, 'h10778, 'h10788, 'h10ab3, 'h10798, 'h10cb8, 'h107a8, 'h10ab4, 'h107b8, 'h107c8, 'h10ab5, 'h107d8, 'h107e8, 'h10ab6, 'h103bc, 'h107f8, 'h10808, 'h10ab7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10818, 'h10828, 'h10ab8, 'h10838, 'h10848, 'h10ab9, 'h10cb8, 'h10858, 'h10868, 'h10aba, 'h10878, 'h10888, 'h10abb, 'h10898, 'h103bc, 'h108a8, 'h10abc, 'h108b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c8, 'h10abd, 'h108d8, 'h106e8, 'h10abe, 'h10cc8, 'h106f8, 'h10708, 'h10abf, 'h10718, 'h10728, 'h10ac0, 'h10738, 'h10748, 'h10ac1, 'h103bc, 'h10758, 'h10768, 'h10ac2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10778, 'h10788, 'h10ac3, 'h10798, 'h10cc8, 'h107a8, 'h10ac4, 'h107b8, 'h107c8, 'h10ac5, 'h107d8, 'h107e8, 'h10ac6, 'h107f8, 'h103bc, 'h10808, 'h10ac7, 'h10818, 'h21f8e, 'h21f8f, 'h21f8d, 'h10828, 'h10ac8, 'h10838, 'h10848, 'h10ac9, 'h10cc8, 'h10858, 'h10868, 'h10aca, 'h10878, 'h10888, 'h10acb, 'h10898, 'h108a8, 'h10acc, 'h103bc, 'h108b8, 'h108c8, 'h10acd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d8, 'h106e8, 'h10ace, 'h10cd8, 'h106f8, 'h10708, 'h10acf, 'h10718, 'h10728, 'h10ad0, 'h10738, 'h10748, 'h10ad1, 'h10758, 'h103bc, 'h10768, 'h10ad2, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10788, 'h10ad3, 'h10798, 'h10cd8, 'h107a8, 'h10ad4, 'h107b8, 'h107c8, 'h10ad5, 'h107d8, 'h107e8, 'h10ad6, 'h107f8, 'h10808, 'h10ad7, 'h103bc, 'h10818, 'h10828, 'h10ad8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10838, 'h10848, 'h10ad9, 'h10cd8, 'h10858, 'h10868, 'h10ada, 'h10878, 'h10888, 'h10adb, 'h10898, 'h108a8, 'h10adc, 'h108b8, 'h103bc, 'h108c8, 'h10add, 'h108d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e9, 'h108de, 'h10ae9, 'h106f9, 'h10709, 'h108df, 'h10719, 'h10729, 'h108e0, 'h10739, 'h10749, 'h108e1, 'h10759, 'h10769, 'h108e2, 'h103bc, 'h10779, 'h10789, 'h108e3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10799, 'h10ae9, 'h107a9, 'h108e4, 'h107b9, 'h107c9, 'h108e5, 'h107d9, 'h107e9, 'h108e6, 'h107f9, 'h10809, 'h108e7, 'h10819, 'h103bc, 'h10829, 'h108e8, 'h10839, 'h21f8e, 'h21f8f, 'h21f8d, 'h10849, 'h108e9, 'h10ae9, 'h10859, 'h10869, 'h108ea, 'h10879, 'h10889, 'h108eb, 'h10899, 'h108a9, 'h108ec, 'h108b9, 'h108c9, 'h108ed, 'h103bc, 'h108d9, 'h106e9, 'h108ee, 'h10af9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f9, 'h10709, 'h108ef, 'h10719, 'h10729, 'h108f0, 'h10739, 'h10749, 'h108f1, 'h10759, 'h10769, 'h108f2, 'h10779, 'h103bc, 'h10789, 'h108f3, 'h10799, 'h10af9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a9, 'h108f4, 'h107b9, 'h107c9, 'h108f5, 'h107d9, 'h107e9, 'h108f6, 'h107f9, 'h10809, 'h108f7, 'h10819, 'h10829, 'h108f8, 'h103bc, 'h10839, 'h10849, 'h108f9, 'h10af9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10859, 'h10869, 'h108fa, 'h10879, 'h10889, 'h108fb, 'h10899, 'h108a9, 'h108fc, 'h108b9, 'h108c9, 'h108fd, 'h108d9, 'h103bc, 'h106e9, 'h108fe, 'h10b09, 'h106f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h108ff, 'h10719, 'h10729, 'h10900, 'h10739, 'h10749, 'h10901, 'h10759, 'h10769, 'h10902, 'h10779, 'h10789, 'h10903, 'h103bc, 'h10799, 'h10b09, 'h107a9, 'h10904, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b9, 'h107c9, 'h10905, 'h107d9, 'h107e9, 'h10906, 'h107f9, 'h10809, 'h10907, 'h10819, 'h10829, 'h10908, 'h10839, 'h103bc, 'h10849, 'h10909, 'h10b09, 'h10859, 'h21f8e, 'h21f8f, 'h21f8d, 'h10869, 'h1090a, 'h10879, 'h10889, 'h1090b, 'h10899, 'h108a9, 'h1090c, 'h108b9, 'h108c9, 'h1090d, 'h108d9, 'h106e9, 'h1090e, 'h10b19, 'h103bc, 'h106f9, 'h10709, 'h1090f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10719, 'h10729, 'h10910, 'h10739, 'h10749, 'h10911, 'h10759, 'h10769, 'h10912, 'h10779, 'h10789, 'h10913, 'h10799, 'h10b19, 'h103bc, 'h107a9, 'h10914, 'h107b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c9, 'h10915, 'h107d9, 'h107e9, 'h10916, 'h107f9, 'h10809, 'h10917, 'h10819, 'h10829, 'h10918, 'h10839, 'h10849, 'h10919, 'h10b19, 'h103bc, 'h10859, 'h10869, 'h1091a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10879, 'h10889, 'h1091b, 'h10899, 'h108a9, 'h1091c, 'h108b9, 'h108c9, 'h1091d, 'h108d9, 'h106e9, 'h1091e, 'h10b29, 'h106f9, 'h103bc, 'h10709, 'h1091f, 'h10719, 'h21f8e, 'h21f8f, 'h21f8d, 'h10729, 'h10920, 'h10739, 'h10749, 'h10921, 'h10759, 'h10769, 'h10922, 'h10779, 'h10789, 'h10923, 'h10799, 'h10b29, 'h107a9, 'h10924, 'h103bc, 'h107b9, 'h107c9, 'h10925, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d9, 'h107e9, 'h10926, 'h107f9, 'h10809, 'h10927, 'h10819, 'h10829, 'h10928, 'h10839, 'h10849, 'h10929, 'h10b29, 'h10859, 'h103bc, 'h10869, 'h1092a, 'h10879, 'h21f8e, 'h21f8f, 'h21f8d, 'h10889, 'h1092b, 'h10899, 'h108a9, 'h1092c, 'h108b9, 'h108c9, 'h1092d, 'h108d9, 'h106e9, 'h1092e, 'h10b39, 'h106f9, 'h10709, 'h1092f, 'h103bc, 'h10719, 'h10729, 'h10930, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10749, 'h10931, 'h10759, 'h10769, 'h10932, 'h10779, 'h10789, 'h10933, 'h10799, 'h10b39, 'h107a9, 'h10934, 'h107b9, 'h103bc, 'h107c9, 'h10935, 'h107d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e9, 'h10936, 'h107f9, 'h10809, 'h10937, 'h10819, 'h10829, 'h10938, 'h10839, 'h10849, 'h10939, 'h10b39, 'h10859, 'h10869, 'h1093a, 'h103bc, 'h10879, 'h10889, 'h1093b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10899, 'h108a9, 'h1093c, 'h108b9, 'h108c9, 'h1093d, 'h108d9, 'h106e9, 'h1093e, 'h10b49, 'h106f9, 'h10709, 'h1093f, 'h10719, 'h103bc, 'h10729, 'h10940, 'h10739, 'h21f8e, 'h21f8f, 'h21f8d, 'h10749, 'h10941, 'h10759, 'h10769, 'h10942, 'h10779, 'h10789, 'h10943, 'h10799, 'h10b49, 'h107a9, 'h10944, 'h107b9, 'h107c9, 'h10945, 'h103bc, 'h107d9, 'h107e9, 'h10946, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f9, 'h10809, 'h10947, 'h10819, 'h10829, 'h10948, 'h10839, 'h10849, 'h10949, 'h10b49, 'h10859, 'h10869, 'h1094a, 'h10879, 'h103bc, 'h10889, 'h1094b, 'h10899, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a9, 'h1094c, 'h108b9, 'h108c9, 'h1094d, 'h108d9, 'h106e9, 'h1094e, 'h10b59, 'h106f9, 'h10709, 'h1094f, 'h10719, 'h10729, 'h10950, 'h103bc, 'h10739, 'h10749, 'h10951, 'h21f8e, 'h21f8f, 'h21f8d, 'h10759, 'h10769, 'h10952, 'h10779, 'h10789, 'h10953, 'h10799, 'h10b59, 'h107a9, 'h10954, 'h107b9, 'h107c9, 'h10955, 'h107d9, 'h103bc, 'h107e9, 'h10956, 'h107f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10809, 'h10957, 'h10819, 'h10829, 'h10958, 'h10839, 'h10849, 'h10959, 'h10b59, 'h10859, 'h10869, 'h1095a, 'h10879, 'h10889, 'h1095b, 'h103bc, 'h10899, 'h108a9, 'h1095c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b9, 'h108c9, 'h1095d, 'h108d9, 'h106e9, 'h1095e, 'h10b69, 'h106f9, 'h10709, 'h1095f, 'h10719, 'h10729, 'h10960, 'h10739, 'h103bc, 'h10749, 'h10961, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h10769, 'h10962, 'h10779, 'h10789, 'h10963, 'h10799, 'h10b69, 'h107a9, 'h10964, 'h107b9, 'h107c9, 'h10965, 'h107d9, 'h107e9, 'h10966, 'h103bc, 'h107f9, 'h10809, 'h10967, 'h21f8e, 'h21f8f, 'h21f8d, 'h10819, 'h10829, 'h10968, 'h10839, 'h10849, 'h10969, 'h10b69, 'h10859, 'h10869, 'h1096a, 'h10879, 'h10889, 'h1096b, 'h10899, 'h103bc, 'h108a9, 'h1096c, 'h108b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c9, 'h1096d, 'h108d9, 'h106e9, 'h1096e, 'h10b79, 'h106f9, 'h10709, 'h1096f, 'h10719, 'h10729, 'h10970, 'h10739, 'h10749, 'h10971, 'h103bc, 'h10759, 'h10769, 'h10972, 'h21f8e, 'h21f8f, 'h21f8d, 'h10779, 'h10789, 'h10973, 'h10799, 'h10b79, 'h107a9, 'h10974, 'h107b9, 'h107c9, 'h10975, 'h107d9, 'h107e9, 'h10976, 'h107f9, 'h103bc, 'h10809, 'h10977, 'h10819, 'h21f8e, 'h21f8f, 'h21f8d, 'h10829, 'h10978, 'h10839, 'h10849, 'h10979, 'h10b79, 'h10859, 'h10869, 'h1097a, 'h10879, 'h10889, 'h1097b, 'h10899, 'h108a9, 'h1097c, 'h103bc, 'h108b9, 'h108c9, 'h1097d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d9, 'h106e9, 'h1097e, 'h10b89, 'h106f9, 'h10709, 'h1097f, 'h10719, 'h10729, 'h10980, 'h10739, 'h10749, 'h10981, 'h10759, 'h103bc, 'h10769, 'h10982, 'h10779, 'h21f8e, 'h21f8f, 'h21f8d, 'h10789, 'h10983, 'h10799, 'h10b89, 'h107a9, 'h10984, 'h107b9, 'h107c9, 'h10985, 'h107d9, 'h107e9, 'h10986, 'h107f9, 'h10809, 'h10987, 'h103bc, 'h10819, 'h10829, 'h10988, 'h21f8e, 'h21f8f, 'h21f8d, 'h10839, 'h10849, 'h10989, 'h10b89, 'h10859, 'h10869, 'h1098a, 'h10879, 'h10889, 'h1098b, 'h10899, 'h108a9, 'h1098c, 'h108b9, 'h103bc, 'h108c9, 'h1098d, 'h108d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e9, 'h1098e, 'h10b99, 'h106f9, 'h10709, 'h1098f, 'h10719, 'h10729, 'h10990, 'h10739, 'h10749, 'h10991, 'h10759, 'h10769, 'h10992, 'h103bc, 'h10779, 'h10789, 'h10993, 'h21f8e, 'h21f8f, 'h21f8d, 'h10799, 'h10b99, 'h107a9, 'h10994, 'h107b9, 'h107c9, 'h10995, 'h107d9, 'h107e9, 'h10996, 'h107f9, 'h10809, 'h10997, 'h10819, 'h103bc, 'h10829, 'h10998, 'h10839, 'h21f8e, 'h21f8f, 'h21f8d, 'h10849, 'h10999, 'h10b99, 'h10859, 'h10869, 'h1099a, 'h10879, 'h10889, 'h1099b, 'h10899, 'h108a9, 'h1099c, 'h108b9, 'h108c9, 'h1099d, 'h103bc, 'h108d9, 'h106e9, 'h1099e, 'h10ba9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f9, 'h10709, 'h1099f, 'h10719, 'h10729, 'h109a0, 'h10739, 'h10749, 'h109a1, 'h10759, 'h10769, 'h109a2, 'h10779, 'h103bc, 'h10789, 'h109a3, 'h10799, 'h10ba9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a9, 'h109a4, 'h107b9, 'h107c9, 'h109a5, 'h107d9, 'h107e9, 'h109a6, 'h107f9, 'h10809, 'h109a7, 'h10819, 'h10829, 'h109a8, 'h103bc, 'h10839, 'h10849, 'h109a9, 'h10ba9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10859, 'h10869, 'h109aa, 'h10879, 'h10889, 'h109ab, 'h10899, 'h108a9, 'h109ac, 'h108b9, 'h108c9, 'h109ad, 'h108d9, 'h103bc, 'h106e9, 'h109ae, 'h10bb9, 'h106f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h109af, 'h10719, 'h10729, 'h109b0, 'h10739, 'h10749, 'h109b1, 'h10759, 'h10769, 'h109b2, 'h10779, 'h10789, 'h109b3, 'h103bc, 'h10799, 'h10bb9, 'h107a9, 'h109b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b9, 'h107c9, 'h109b5, 'h107d9, 'h107e9, 'h109b6, 'h107f9, 'h10809, 'h109b7, 'h10819, 'h10829, 'h109b8, 'h10839, 'h103bc, 'h10849, 'h109b9, 'h10bb9, 'h10859, 'h21f8e, 'h21f8f, 'h21f8d, 'h10869, 'h109ba, 'h10879, 'h10889, 'h109bb, 'h10899, 'h108a9, 'h109bc, 'h108b9, 'h108c9, 'h109bd, 'h108d9, 'h106e9, 'h109be, 'h10bc9, 'h103bc, 'h106f9, 'h10709, 'h109bf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10719, 'h10729, 'h109c0, 'h10739, 'h10749, 'h109c1, 'h10759, 'h10769, 'h109c2, 'h10779, 'h10789, 'h109c3, 'h10799, 'h10bc9, 'h103bc, 'h107a9, 'h109c4, 'h107b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c9, 'h109c5, 'h107d9, 'h107e9, 'h109c6, 'h107f9, 'h10809, 'h109c7, 'h10819, 'h10829, 'h109c8, 'h10839, 'h10849, 'h109c9, 'h10bc9, 'h103bc, 'h10859, 'h10869, 'h109ca, 'h21f8e, 'h21f8f, 'h21f8d, 'h10879, 'h10889, 'h109cb, 'h10899, 'h108a9, 'h109cc, 'h108b9, 'h108c9, 'h109cd, 'h108d9, 'h106e9, 'h109ce, 'h10bd9, 'h106f9, 'h103bc, 'h10709, 'h109cf, 'h10719, 'h21f8e, 'h21f8f, 'h21f8d, 'h10729, 'h109d0, 'h10739, 'h10749, 'h109d1, 'h10759, 'h10769, 'h109d2, 'h10779, 'h10789, 'h109d3, 'h10799, 'h10bd9, 'h107a9, 'h109d4, 'h103bc, 'h107b9, 'h107c9, 'h109d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d9, 'h107e9, 'h109d6, 'h107f9, 'h10809, 'h109d7, 'h10819, 'h10829, 'h109d8, 'h10839, 'h10849, 'h109d9, 'h10bd9, 'h10859, 'h103bc, 'h10869, 'h109da, 'h10879, 'h21f8e, 'h21f8f, 'h21f8d, 'h10889, 'h109db, 'h10899, 'h108a9, 'h109dc, 'h108b9, 'h108c9, 'h109dd, 'h108d9, 'h106e9, 'h109de, 'h10be9, 'h106f9, 'h10709, 'h109df, 'h103bc, 'h10719, 'h10729, 'h109e0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10749, 'h109e1, 'h10759, 'h10769, 'h109e2, 'h10779, 'h10789, 'h109e3, 'h10799, 'h10be9, 'h107a9, 'h109e4, 'h107b9, 'h103bc, 'h107c9, 'h109e5, 'h107d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e9, 'h109e6, 'h107f9, 'h10809, 'h109e7, 'h10819, 'h10829, 'h109e8, 'h10839, 'h10849, 'h109e9, 'h10be9, 'h10859, 'h10869, 'h109ea, 'h103bc, 'h10879, 'h10889, 'h109eb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10899, 'h108a9, 'h109ec, 'h108b9, 'h108c9, 'h109ed, 'h108d9, 'h106e9, 'h109ee, 'h10bf9, 'h106f9, 'h10709, 'h109ef, 'h10719, 'h103bc, 'h10729, 'h109f0, 'h10739, 'h21f8e, 'h21f8f, 'h21f8d, 'h10749, 'h109f1, 'h10759, 'h10769, 'h109f2, 'h10779, 'h10789, 'h109f3, 'h10799, 'h10bf9, 'h107a9, 'h109f4, 'h107b9, 'h107c9, 'h109f5, 'h103bc, 'h107d9, 'h107e9, 'h109f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f9, 'h10809, 'h109f7, 'h10819, 'h10829, 'h109f8, 'h10839, 'h10849, 'h109f9, 'h10bf9, 'h10859, 'h10869, 'h109fa, 'h10879, 'h103bc, 'h10889, 'h109fb, 'h10899, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a9, 'h109fc, 'h108b9, 'h108c9, 'h109fd, 'h108d9, 'h106e9, 'h109fe, 'h10c09, 'h106f9, 'h10709, 'h109ff, 'h10719, 'h10729, 'h10a00, 'h103bc, 'h10739, 'h10749, 'h10a01, 'h21f8e, 'h21f8f, 'h21f8d, 'h10759, 'h10769, 'h10a02, 'h10779, 'h10789, 'h10a03, 'h10799, 'h10c09, 'h107a9, 'h10a04, 'h107b9, 'h107c9, 'h10a05, 'h107d9, 'h103bc, 'h107e9, 'h10a06, 'h107f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10809, 'h10a07, 'h10819, 'h10829, 'h10a08, 'h10839, 'h10849, 'h10a09, 'h10c09, 'h10859, 'h10869, 'h10a0a, 'h10879, 'h10889, 'h10a0b, 'h103bc, 'h10899, 'h108a9, 'h10a0c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b9, 'h108c9, 'h10a0d, 'h108d9, 'h106e9, 'h10a0e, 'h10c19, 'h106f9, 'h10709, 'h10a0f, 'h10719, 'h10729, 'h10a10, 'h10739, 'h103bc, 'h10749, 'h10a11, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h10769, 'h10a12, 'h10779, 'h10789, 'h10a13, 'h10799, 'h10c19, 'h107a9, 'h10a14, 'h107b9, 'h107c9, 'h10a15, 'h107d9, 'h107e9, 'h10a16, 'h103bc, 'h107f9, 'h10809, 'h10a17, 'h21f8e, 'h21f8f, 'h21f8d, 'h10819, 'h10829, 'h10a18, 'h10839, 'h10849, 'h10a19, 'h10c19, 'h10859, 'h10869, 'h10a1a, 'h10879, 'h10889, 'h10a1b, 'h10899, 'h103bc, 'h108a9, 'h10a1c, 'h108b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c9, 'h10a1d, 'h108d9, 'h106e9, 'h10a1e, 'h10c29, 'h106f9, 'h10709, 'h10a1f, 'h10719, 'h10729, 'h10a20, 'h10739, 'h10749, 'h10a21, 'h103bc, 'h10759, 'h10769, 'h10a22, 'h21f8e, 'h21f8f, 'h21f8d, 'h10779, 'h10789, 'h10a23, 'h10799, 'h10c29, 'h107a9, 'h10a24, 'h107b9, 'h107c9, 'h10a25, 'h107d9, 'h107e9, 'h10a26, 'h107f9, 'h103bc, 'h10809, 'h10a27, 'h10819, 'h21f8e, 'h21f8f, 'h21f8d, 'h10829, 'h10a28, 'h10839, 'h10849, 'h10a29, 'h10c29, 'h10859, 'h10869, 'h10a2a, 'h10879, 'h10889, 'h10a2b, 'h10899, 'h108a9, 'h10a2c, 'h103bc, 'h108b9, 'h108c9, 'h10a2d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d9, 'h106e9, 'h10a2e, 'h10c39, 'h106f9, 'h10709, 'h10a2f, 'h10719, 'h10729, 'h10a30, 'h10739, 'h10749, 'h10a31, 'h10759, 'h103bc, 'h10769, 'h10a32, 'h10779, 'h21f8e, 'h21f8f, 'h21f8d, 'h10789, 'h10a33, 'h10799, 'h10c39, 'h107a9, 'h10a34, 'h107b9, 'h107c9, 'h10a35, 'h107d9, 'h107e9, 'h10a36, 'h107f9, 'h10809, 'h10a37, 'h103bc, 'h10819, 'h10829, 'h10a38, 'h21f8e, 'h21f8f, 'h21f8d, 'h10839, 'h10849, 'h10a39, 'h10c39, 'h10859, 'h10869, 'h10a3a, 'h10879, 'h10889, 'h10a3b, 'h10899, 'h108a9, 'h10a3c, 'h108b9, 'h103bc, 'h108c9, 'h10a3d, 'h108d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e9, 'h10a3e, 'h10c49, 'h106f9, 'h10709, 'h10a3f, 'h10719, 'h10729, 'h10a40, 'h10739, 'h10749, 'h10a41, 'h10759, 'h10769, 'h10a42, 'h103bc, 'h10779, 'h10789, 'h10a43, 'h21f8e, 'h21f8f, 'h21f8d, 'h10799, 'h10c49, 'h107a9, 'h10a44, 'h107b9, 'h107c9, 'h10a45, 'h107d9, 'h107e9, 'h10a46, 'h107f9, 'h10809, 'h10a47, 'h10819, 'h103bc, 'h10829, 'h10a48, 'h10839, 'h21f8e, 'h21f8f, 'h21f8d, 'h10849, 'h10a49, 'h10c49, 'h10859, 'h10869, 'h10a4a, 'h10879, 'h10889, 'h10a4b, 'h10899, 'h108a9, 'h10a4c, 'h108b9, 'h108c9, 'h10a4d, 'h103bc, 'h108d9, 'h106e9, 'h10a4e, 'h10c59, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f9, 'h10709, 'h10a4f, 'h10719, 'h10729, 'h10a50, 'h10739, 'h10749, 'h10a51, 'h10759, 'h10769, 'h10a52, 'h10779, 'h103bc, 'h10789, 'h10a53, 'h10799, 'h10c59, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a9, 'h10a54, 'h107b9, 'h107c9, 'h10a55, 'h107d9, 'h107e9, 'h10a56, 'h107f9, 'h10809, 'h10a57, 'h10819, 'h10829, 'h10a58, 'h103bc, 'h10839, 'h10849, 'h10a59, 'h10c59, 'h21f8e, 'h21f8f, 'h21f8d, 'h10859, 'h10869, 'h10a5a, 'h10879, 'h10889, 'h10a5b, 'h10899, 'h108a9, 'h10a5c, 'h108b9, 'h108c9, 'h10a5d, 'h108d9, 'h103bc, 'h106e9, 'h10a5e, 'h10c69, 'h106f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10a5f, 'h10719, 'h10729, 'h10a60, 'h10739, 'h10749, 'h10a61, 'h10759, 'h10769, 'h10a62, 'h10779, 'h10789, 'h10a63, 'h103bc, 'h10799, 'h10c69, 'h107a9, 'h10a64, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b9, 'h107c9, 'h10a65, 'h107d9, 'h107e9, 'h10a66, 'h107f9, 'h10809, 'h10a67, 'h10819, 'h10829, 'h10a68, 'h10839, 'h103bc, 'h10849, 'h10a69, 'h10c69, 'h10859, 'h21f8e, 'h21f8f, 'h21f8d, 'h10869, 'h10a6a, 'h10879, 'h10889, 'h10a6b, 'h10899, 'h108a9, 'h10a6c, 'h108b9, 'h108c9, 'h10a6d, 'h108d9, 'h106e9, 'h10a6e, 'h10c79, 'h103bc, 'h106f9, 'h10709, 'h10a6f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10719, 'h10729, 'h10a70, 'h10739, 'h10749, 'h10a71, 'h10759, 'h10769, 'h10a72, 'h10779, 'h10789, 'h10a73, 'h10799, 'h10c79, 'h103bc, 'h107a9, 'h10a74, 'h107b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c9, 'h10a75, 'h107d9, 'h107e9, 'h10a76, 'h107f9, 'h10809, 'h10a77, 'h10819, 'h10829, 'h10a78, 'h10839, 'h10849, 'h10a79, 'h10c79, 'h103bc, 'h10859, 'h10869, 'h10a7a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10879, 'h10889, 'h10a7b, 'h10899, 'h108a9, 'h10a7c, 'h108b9, 'h108c9, 'h10a7d, 'h108d9, 'h106e9, 'h10a7e, 'h10c89, 'h106f9, 'h103bc, 'h10709, 'h10a7f, 'h10719, 'h21f8e, 'h21f8f, 'h21f8d, 'h10729, 'h10a80, 'h10739, 'h10749, 'h10a81, 'h10759, 'h10769, 'h10a82, 'h10779, 'h10789, 'h10a83, 'h10799, 'h10c89, 'h107a9, 'h10a84, 'h103bc, 'h107b9, 'h107c9, 'h10a85, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d9, 'h107e9, 'h10a86, 'h107f9, 'h10809, 'h10a87, 'h10819, 'h10829, 'h10a88, 'h10839, 'h10849, 'h10a89, 'h10c89, 'h10859, 'h103bc, 'h10869, 'h10a8a, 'h10879, 'h21f8e, 'h21f8f, 'h21f8d, 'h10889, 'h10a8b, 'h10899, 'h108a9, 'h10a8c, 'h108b9, 'h108c9, 'h10a8d, 'h108d9, 'h106e9, 'h10a8e, 'h10c99, 'h106f9, 'h10709, 'h10a8f, 'h103bc, 'h10719, 'h10729, 'h10a90, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10749, 'h10a91, 'h10759, 'h10769, 'h10a92, 'h10779, 'h10789, 'h10a93, 'h10799, 'h10c99, 'h107a9, 'h10a94, 'h107b9, 'h103bc, 'h107c9, 'h10a95, 'h107d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e9, 'h10a96, 'h107f9, 'h10809, 'h10a97, 'h10819, 'h10829, 'h10a98, 'h10839, 'h10849, 'h10a99, 'h10c99, 'h10859, 'h10869, 'h10a9a, 'h103bc, 'h10879, 'h10889, 'h10a9b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10899, 'h108a9, 'h10a9c, 'h108b9, 'h108c9, 'h10a9d, 'h108d9, 'h106e9, 'h10a9e, 'h10ca9, 'h106f9, 'h10709, 'h10a9f, 'h10719, 'h103bc, 'h10729, 'h10aa0, 'h10739, 'h21f8e, 'h21f8f, 'h21f8d, 'h10749, 'h10aa1, 'h10759, 'h10769, 'h10aa2, 'h10779, 'h10789, 'h10aa3, 'h10799, 'h10ca9, 'h107a9, 'h10aa4, 'h107b9, 'h107c9, 'h10aa5, 'h103bc, 'h107d9, 'h107e9, 'h10aa6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f9, 'h10809, 'h10aa7, 'h10819, 'h10829, 'h10aa8, 'h10839, 'h10849, 'h10aa9, 'h10ca9, 'h10859, 'h10869, 'h10aaa, 'h10879, 'h103bc, 'h10889, 'h10aab, 'h10899, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a9, 'h10aac, 'h108b9, 'h108c9, 'h10aad, 'h108d9, 'h106e9, 'h10aae, 'h10cb9, 'h106f9, 'h10709, 'h10aaf, 'h10719, 'h10729, 'h10ab0, 'h103bc, 'h10739, 'h10749, 'h10ab1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10759, 'h10769, 'h10ab2, 'h10779, 'h10789, 'h10ab3, 'h10799, 'h10cb9, 'h107a9, 'h10ab4, 'h107b9, 'h107c9, 'h10ab5, 'h107d9, 'h103bc, 'h107e9, 'h10ab6, 'h107f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10809, 'h10ab7, 'h10819, 'h10829, 'h10ab8, 'h10839, 'h10849, 'h10ab9, 'h10cb9, 'h10859, 'h10869, 'h10aba, 'h10879, 'h10889, 'h10abb, 'h103bc, 'h10899, 'h108a9, 'h10abc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b9, 'h108c9, 'h10abd, 'h108d9, 'h106e9, 'h10abe, 'h10cc9, 'h106f9, 'h10709, 'h10abf, 'h10719, 'h10729, 'h10ac0, 'h10739, 'h103bc, 'h10749, 'h10ac1, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h10769, 'h10ac2, 'h10779, 'h10789, 'h10ac3, 'h10799, 'h10cc9, 'h107a9, 'h10ac4, 'h107b9, 'h107c9, 'h10ac5, 'h107d9, 'h107e9, 'h10ac6, 'h103bc, 'h107f9, 'h10809, 'h10ac7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10819, 'h10829, 'h10ac8, 'h10839, 'h10849, 'h10ac9, 'h10cc9, 'h10859, 'h10869, 'h10aca, 'h10879, 'h10889, 'h10acb, 'h10899, 'h103bc, 'h108a9, 'h10acc, 'h108b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c9, 'h10acd, 'h108d9, 'h106e9, 'h10ace, 'h10cd9, 'h106f9, 'h10709, 'h10acf, 'h10719, 'h10729, 'h10ad0, 'h10739, 'h10749, 'h10ad1, 'h103bc, 'h10759, 'h10769, 'h10ad2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10779, 'h10789, 'h10ad3, 'h10799, 'h10cd9, 'h107a9, 'h10ad4, 'h107b9, 'h107c9, 'h10ad5, 'h107d9, 'h107e9, 'h10ad6, 'h107f9, 'h103bc, 'h10809, 'h10ad7, 'h10819, 'h21f8e, 'h21f8f, 'h21f8d, 'h10829, 'h10ad8, 'h10839, 'h10849, 'h10ad9, 'h10cd9, 'h10859, 'h10869, 'h10ada, 'h10879, 'h10889, 'h10adb, 'h10899, 'h108a9, 'h10adc, 'h103bc, 'h108b9, 'h108c9, 'h10add, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d9, 'h106e9, 'h108de, 'h10ae9, 'h106f9, 'h10709, 'h108df, 'h10719, 'h10729, 'h108e0, 'h10739, 'h10749, 'h108e1, 'h10759, 'h103bc, 'h10769, 'h108e2, 'h10779, 'h21f8e, 'h21f8f, 'h21f8d, 'h10789, 'h108e3, 'h10799, 'h10ae9, 'h107a9, 'h108e4, 'h107b9, 'h107c9, 'h108e5, 'h107d9, 'h107e9, 'h108e6, 'h107f9, 'h10809, 'h108e7, 'h103bc, 'h10819, 'h10829, 'h108e8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10839, 'h10849, 'h108e9, 'h10ae9, 'h10859, 'h10869, 'h108ea, 'h10879, 'h10889, 'h108eb, 'h10899, 'h108a9, 'h108ec, 'h108b9, 'h103bc, 'h108c9, 'h108ed, 'h108d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e9, 'h108ee, 'h10af9, 'h106f9, 'h10709, 'h108ef, 'h10719, 'h10729, 'h108f0, 'h10739, 'h10749, 'h108f1, 'h10759, 'h10769, 'h108f2, 'h103bc, 'h10779, 'h10789, 'h108f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10799, 'h10af9, 'h107a9, 'h108f4, 'h107b9, 'h107c9, 'h108f5, 'h107d9, 'h107e9, 'h108f6, 'h107f9, 'h10809, 'h108f7, 'h10819, 'h103bc, 'h10829, 'h108f8, 'h10839, 'h21f8e, 'h21f8f, 'h21f8d, 'h10849, 'h108f9, 'h10af9, 'h10859, 'h10869, 'h108fa, 'h10879, 'h10889, 'h108fb, 'h10899, 'h108a9, 'h108fc, 'h108b9, 'h108c9, 'h108fd, 'h103bc, 'h108d9, 'h106e9, 'h108fe, 'h10b09, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f9, 'h10709, 'h108ff, 'h10719, 'h10729, 'h10900, 'h10739, 'h10749, 'h10901, 'h10759, 'h10769, 'h10902, 'h10779, 'h103bc, 'h10789, 'h10903, 'h10799, 'h10b09, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a9, 'h10904, 'h107b9, 'h107c9, 'h10905, 'h107d9, 'h107e9, 'h10906, 'h107f9, 'h10809, 'h10907, 'h10819, 'h10829, 'h10908, 'h103bc, 'h10839, 'h10849, 'h10909, 'h10b09, 'h21f8e, 'h21f8f, 'h21f8d, 'h10859, 'h10869, 'h1090a, 'h10879, 'h10889, 'h1090b, 'h10899, 'h108a9, 'h1090c, 'h108b9, 'h108c9, 'h1090d, 'h108d9, 'h103bc, 'h106e9, 'h1090e, 'h10b19, 'h106f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h1090f, 'h10719, 'h10729, 'h10910, 'h10739, 'h10749, 'h10911, 'h10759, 'h10769, 'h10912, 'h10779, 'h10789, 'h10913, 'h103bc, 'h10799, 'h10b19, 'h107a9, 'h10914, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b9, 'h107c9, 'h10915, 'h107d9, 'h107e9, 'h10916, 'h107f9, 'h10809, 'h10917, 'h10819, 'h10829, 'h10918, 'h10839, 'h103bc, 'h10849, 'h10919, 'h10b19, 'h10859, 'h21f8e, 'h21f8f, 'h21f8d, 'h10869, 'h1091a, 'h10879, 'h10889, 'h1091b, 'h10899, 'h108a9, 'h1091c, 'h108b9, 'h108c9, 'h1091d, 'h108d9, 'h106e9, 'h1091e, 'h10b29, 'h103bc, 'h106f9, 'h10709, 'h1091f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10719, 'h10729, 'h10920, 'h10739, 'h10749, 'h10921, 'h10759, 'h10769, 'h10922, 'h10779, 'h10789, 'h10923, 'h10799, 'h10b29, 'h103bc, 'h107a9, 'h10924, 'h107b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c9, 'h10925, 'h107d9, 'h107e9, 'h10926, 'h107f9, 'h10809, 'h10927, 'h10819, 'h10829, 'h10928, 'h10839, 'h10849, 'h10929, 'h10b29, 'h103bc, 'h10859, 'h10869, 'h1092a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10879, 'h10889, 'h1092b, 'h10899, 'h108a9, 'h1092c, 'h108b9, 'h108c9, 'h1092d, 'h108d9, 'h106e9, 'h1092e, 'h10b39, 'h106f9, 'h103bc, 'h10709, 'h1092f, 'h10719, 'h21f8e, 'h21f8f, 'h21f8d, 'h10729, 'h10930, 'h10739, 'h10749, 'h10931, 'h10759, 'h10769, 'h10932, 'h10779, 'h10789, 'h10933, 'h10799, 'h10b39, 'h107a9, 'h10934, 'h103bc, 'h107b9, 'h107c9, 'h10935, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d9, 'h107e9, 'h10936, 'h107f9, 'h10809, 'h10937, 'h10819, 'h10829, 'h10938, 'h10839, 'h10849, 'h10939, 'h10b39, 'h10859, 'h103bc, 'h10869, 'h1093a, 'h10879, 'h21f8e, 'h21f8f, 'h21f8d, 'h10889, 'h1093b, 'h10899, 'h108a9, 'h1093c, 'h108b9, 'h108c9, 'h1093d, 'h108d9, 'h106e9, 'h1093e, 'h10b49, 'h106f9, 'h10709, 'h1093f, 'h103bc, 'h10719, 'h10729, 'h10940, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10749, 'h10941, 'h10759, 'h10769, 'h10942, 'h10779, 'h10789, 'h10943, 'h10799, 'h10b49, 'h107a9, 'h10944, 'h107b9, 'h103bc, 'h107c9, 'h10945, 'h107d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e9, 'h10946, 'h107f9, 'h10809, 'h10947, 'h10819, 'h10829, 'h10948, 'h10839, 'h10849, 'h10949, 'h10b49, 'h10859, 'h10869, 'h1094a, 'h103bc, 'h10879, 'h10889, 'h1094b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10899, 'h108a9, 'h1094c, 'h108b9, 'h108c9, 'h1094d, 'h108d9, 'h106e9, 'h1094e, 'h10b59, 'h106f9, 'h10709, 'h1094f, 'h10719, 'h103bc, 'h10729, 'h10950, 'h10739, 'h21f8e, 'h21f8f, 'h21f8d, 'h10749, 'h10951, 'h10759, 'h10769, 'h10952, 'h10779, 'h10789, 'h10953, 'h10799, 'h10b59, 'h107a9, 'h10954, 'h107b9, 'h107c9, 'h10955, 'h103bc, 'h107d9, 'h107e9, 'h10956, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f9, 'h10809, 'h10957, 'h10819, 'h10829, 'h10958, 'h10839, 'h10849, 'h10959, 'h10b59, 'h10859, 'h10869, 'h1095a, 'h10879, 'h103bc, 'h10889, 'h1095b, 'h10899, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a9, 'h1095c, 'h108b9, 'h108c9, 'h1095d, 'h108d9, 'h106e9, 'h1095e, 'h10b69, 'h106f9, 'h10709, 'h1095f, 'h10719, 'h10729, 'h10960, 'h103bc, 'h10739, 'h10749, 'h10961, 'h21f8e, 'h21f8f, 'h21f8d, 'h10759, 'h10769, 'h10962, 'h10779, 'h10789, 'h10963, 'h10799, 'h10b69, 'h107a9, 'h10964, 'h107b9, 'h107c9, 'h10965, 'h107d9, 'h103bc, 'h107e9, 'h10966, 'h107f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10809, 'h10967, 'h10819, 'h10829, 'h10968, 'h10839, 'h10849, 'h10969, 'h10b69, 'h10859, 'h10869, 'h1096a, 'h10879, 'h10889, 'h1096b, 'h103bc, 'h10899, 'h108a9, 'h1096c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b9, 'h108c9, 'h1096d, 'h108d9, 'h106e9, 'h1096e, 'h10b79, 'h106f9, 'h10709, 'h1096f, 'h10719, 'h10729, 'h10970, 'h10739, 'h103bc, 'h10749, 'h10971, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h10769, 'h10972, 'h10779, 'h10789, 'h10973, 'h10799, 'h10b79, 'h107a9, 'h10974, 'h107b9, 'h107c9, 'h10975, 'h107d9, 'h107e9, 'h10976, 'h103bc, 'h107f9, 'h10809, 'h10977, 'h21f8e, 'h21f8f, 'h21f8d, 'h10819, 'h10829, 'h10978, 'h10839, 'h10849, 'h10979, 'h10b79, 'h10859, 'h10869, 'h1097a, 'h10879, 'h10889, 'h1097b, 'h10899, 'h103bc, 'h108a9, 'h1097c, 'h108b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c9, 'h1097d, 'h108d9, 'h106e9, 'h1097e, 'h10b89, 'h106f9, 'h10709, 'h1097f, 'h10719, 'h10729, 'h10980, 'h10739, 'h10749, 'h10981, 'h103bc, 'h10759, 'h10769, 'h10982, 'h21f8e, 'h21f8f, 'h21f8d, 'h10779, 'h10789, 'h10983, 'h10799, 'h10b89, 'h107a9, 'h10984, 'h107b9, 'h107c9, 'h10985, 'h107d9, 'h107e9, 'h10986, 'h107f9, 'h103bc, 'h10809, 'h10987, 'h10819, 'h21f8e, 'h21f8f, 'h21f8d, 'h10829, 'h10988, 'h10839, 'h10849, 'h10989, 'h10b89, 'h10859, 'h10869, 'h1098a, 'h10879, 'h10889, 'h1098b, 'h10899, 'h108a9, 'h1098c, 'h103bc, 'h108b9, 'h108c9, 'h1098d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d9, 'h106e9, 'h1098e, 'h10b99, 'h106f9, 'h10709, 'h1098f, 'h10719, 'h10729, 'h10990, 'h10739, 'h10749, 'h10991, 'h10759, 'h103bc, 'h10769, 'h10992, 'h10779, 'h21f8e, 'h21f8f, 'h21f8d, 'h10789, 'h10993, 'h10799, 'h10b99, 'h107a9, 'h10994, 'h107b9, 'h107c9, 'h10995, 'h107d9, 'h107e9, 'h10996, 'h107f9, 'h10809, 'h10997, 'h103bc, 'h10819, 'h10829, 'h10998, 'h21f8e, 'h21f8f, 'h21f8d, 'h10839, 'h10849, 'h10999, 'h10b99, 'h10859, 'h10869, 'h1099a, 'h10879, 'h10889, 'h1099b, 'h10899, 'h108a9, 'h1099c, 'h108b9, 'h103bc, 'h108c9, 'h1099d, 'h108d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e9, 'h1099e, 'h10ba9, 'h106f9, 'h10709, 'h1099f, 'h10719, 'h10729, 'h109a0, 'h10739, 'h10749, 'h109a1, 'h10759, 'h10769, 'h109a2, 'h103bc, 'h10779, 'h10789, 'h109a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10799, 'h10ba9, 'h107a9, 'h109a4, 'h107b9, 'h107c9, 'h109a5, 'h107d9, 'h107e9, 'h109a6, 'h107f9, 'h10809, 'h109a7, 'h10819, 'h103bc, 'h10829, 'h109a8, 'h10839, 'h21f8e, 'h21f8f, 'h21f8d, 'h10849, 'h109a9, 'h10ba9, 'h10859, 'h10869, 'h109aa, 'h10879, 'h10889, 'h109ab, 'h10899, 'h108a9, 'h109ac, 'h108b9, 'h108c9, 'h109ad, 'h103bc, 'h108d9, 'h106e9, 'h109ae, 'h10bb9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f9, 'h10709, 'h109af, 'h10719, 'h10729, 'h109b0, 'h10739, 'h10749, 'h109b1, 'h10759, 'h10769, 'h109b2, 'h10779, 'h103bc, 'h10789, 'h109b3, 'h10799, 'h10bb9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a9, 'h109b4, 'h107b9, 'h107c9, 'h109b5, 'h107d9, 'h107e9, 'h109b6, 'h107f9, 'h10809, 'h109b7, 'h10819, 'h10829, 'h109b8, 'h103bc, 'h10839, 'h10849, 'h109b9, 'h10bb9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10859, 'h10869, 'h109ba, 'h10879, 'h10889, 'h109bb, 'h10899, 'h108a9, 'h109bc, 'h108b9, 'h108c9, 'h109bd, 'h108d9, 'h103bc, 'h106e9, 'h109be, 'h10bc9, 'h106f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h109bf, 'h10719, 'h10729, 'h109c0, 'h10739, 'h10749, 'h109c1, 'h10759, 'h10769, 'h109c2, 'h10779, 'h10789, 'h109c3, 'h103bc, 'h10799, 'h10bc9, 'h107a9, 'h109c4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b9, 'h107c9, 'h109c5, 'h107d9, 'h107e9, 'h109c6, 'h107f9, 'h10809, 'h109c7, 'h10819, 'h10829, 'h109c8, 'h10839, 'h103bc, 'h10849, 'h109c9, 'h10bc9, 'h10859, 'h21f8e, 'h21f8f, 'h21f8d, 'h10869, 'h109ca, 'h10879, 'h10889, 'h109cb, 'h10899, 'h108a9, 'h109cc, 'h108b9, 'h108c9, 'h109cd, 'h108d9, 'h106e9, 'h109ce, 'h10bd9, 'h103bc, 'h106f9, 'h10709, 'h109cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10719, 'h10729, 'h109d0, 'h10739, 'h10749, 'h109d1, 'h10759, 'h10769, 'h109d2, 'h10779, 'h10789, 'h109d3, 'h10799, 'h10bd9, 'h103bc, 'h107a9, 'h109d4, 'h107b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c9, 'h109d5, 'h107d9, 'h107e9, 'h109d6, 'h107f9, 'h10809, 'h109d7, 'h10819, 'h10829, 'h109d8, 'h10839, 'h10849, 'h109d9, 'h10bd9, 'h103bc, 'h10859, 'h10869, 'h109da, 'h21f8e, 'h21f8f, 'h21f8d, 'h10879, 'h10889, 'h109db, 'h10899, 'h108a9, 'h109dc, 'h108b9, 'h108c9, 'h109dd, 'h108d9, 'h106e9, 'h109de, 'h10be9, 'h106f9, 'h103bc, 'h10709, 'h109df, 'h10719, 'h21f8e, 'h21f8f, 'h21f8d, 'h10729, 'h109e0, 'h10739, 'h10749, 'h109e1, 'h10759, 'h10769, 'h109e2, 'h10779, 'h10789, 'h109e3, 'h10799, 'h10be9, 'h107a9, 'h109e4, 'h103bc, 'h107b9, 'h107c9, 'h109e5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d9, 'h107e9, 'h109e6, 'h107f9, 'h10809, 'h109e7, 'h10819, 'h10829, 'h109e8, 'h10839, 'h10849, 'h109e9, 'h10be9, 'h10859, 'h103bc, 'h10869, 'h109ea, 'h10879, 'h21f8e, 'h21f8f, 'h21f8d, 'h10889, 'h109eb, 'h10899, 'h108a9, 'h109ec, 'h108b9, 'h108c9, 'h109ed, 'h108d9, 'h106e9, 'h109ee, 'h10bf9, 'h106f9, 'h10709, 'h109ef, 'h103bc, 'h10719, 'h10729, 'h109f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10749, 'h109f1, 'h10759, 'h10769, 'h109f2, 'h10779, 'h10789, 'h109f3, 'h10799, 'h10bf9, 'h107a9, 'h109f4, 'h107b9, 'h103bc, 'h107c9, 'h109f5, 'h107d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e9, 'h109f6, 'h107f9, 'h10809, 'h109f7, 'h10819, 'h10829, 'h109f8, 'h10839, 'h10849, 'h109f9, 'h10bf9, 'h10859, 'h10869, 'h109fa, 'h103bc, 'h10879, 'h10889, 'h109fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10899, 'h108a9, 'h109fc, 'h108b9, 'h108c9, 'h109fd, 'h108d9, 'h106e9, 'h109fe, 'h10c09, 'h106f9, 'h10709, 'h109ff, 'h10719, 'h103bc, 'h10729, 'h10a00, 'h10739, 'h21f8e, 'h21f8f, 'h21f8d, 'h10749, 'h10a01, 'h10759, 'h10769, 'h10a02, 'h10779, 'h10789, 'h10a03, 'h10799, 'h10c09, 'h107a9, 'h10a04, 'h107b9, 'h107c9, 'h10a05, 'h103bc, 'h107d9, 'h107e9, 'h10a06, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f9, 'h10809, 'h10a07, 'h10819, 'h10829, 'h10a08, 'h10839, 'h10849, 'h10a09, 'h10c09, 'h10859, 'h10869, 'h10a0a, 'h10879, 'h103bc, 'h10889, 'h10a0b, 'h10899, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a9, 'h10a0c, 'h108b9, 'h108c9, 'h10a0d, 'h108d9, 'h106e9, 'h10a0e, 'h10c19, 'h106f9, 'h10709, 'h10a0f, 'h10719, 'h10729, 'h10a10, 'h103bc, 'h10739, 'h10749, 'h10a11, 'h21f8e, 'h21f8f, 'h21f8d, 'h10759, 'h10769, 'h10a12, 'h10779, 'h10789, 'h10a13, 'h10799, 'h10c19, 'h107a9, 'h10a14, 'h107b9, 'h107c9, 'h10a15, 'h107d9, 'h103bc, 'h107e9, 'h10a16, 'h107f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10809, 'h10a17, 'h10819, 'h10829, 'h10a18, 'h10839, 'h10849, 'h10a19, 'h10c19, 'h10859, 'h10869, 'h10a1a, 'h10879, 'h10889, 'h10a1b, 'h103bc, 'h10899, 'h108a9, 'h10a1c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b9, 'h108c9, 'h10a1d, 'h108d9, 'h106e9, 'h10a1e, 'h10c29, 'h106f9, 'h10709, 'h10a1f, 'h10719, 'h10729, 'h10a20, 'h10739, 'h103bc, 'h10749, 'h10a21, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h10769, 'h10a22, 'h10779, 'h10789, 'h10a23, 'h10799, 'h10c29, 'h107a9, 'h10a24, 'h107b9, 'h107c9, 'h10a25, 'h107d9, 'h107e9, 'h10a26, 'h103bc, 'h107f9, 'h10809, 'h10a27, 'h21f8e, 'h21f8f, 'h21f8d, 'h10819, 'h10829, 'h10a28, 'h10839, 'h10849, 'h10a29, 'h10c29, 'h10859, 'h10869, 'h10a2a, 'h10879, 'h10889, 'h10a2b, 'h10899, 'h103bc, 'h108a9, 'h10a2c, 'h108b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c9, 'h10a2d, 'h108d9, 'h106e9, 'h10a2e, 'h10c39, 'h106f9, 'h10709, 'h10a2f, 'h10719, 'h10729, 'h10a30, 'h10739, 'h10749, 'h10a31, 'h103bc, 'h10759, 'h10769, 'h10a32, 'h21f8e, 'h21f8f, 'h21f8d, 'h10779, 'h10789, 'h10a33, 'h10799, 'h10c39, 'h107a9, 'h10a34, 'h107b9, 'h107c9, 'h10a35, 'h107d9, 'h107e9, 'h10a36, 'h107f9, 'h103bc, 'h10809, 'h10a37, 'h10819, 'h21f8e, 'h21f8f, 'h21f8d, 'h10829, 'h10a38, 'h10839, 'h10849, 'h10a39, 'h10c39, 'h10859, 'h10869, 'h10a3a, 'h10879, 'h10889, 'h10a3b, 'h10899, 'h108a9, 'h10a3c, 'h103bc, 'h108b9, 'h108c9, 'h10a3d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d9, 'h106e9, 'h10a3e, 'h10c49, 'h106f9, 'h10709, 'h10a3f, 'h10719, 'h10729, 'h10a40, 'h10739, 'h10749, 'h10a41, 'h10759, 'h103bc, 'h10769, 'h10a42, 'h10779, 'h21f8e, 'h21f8f, 'h21f8d, 'h10789, 'h10a43, 'h10799, 'h10c49, 'h107a9, 'h10a44, 'h107b9, 'h107c9, 'h10a45, 'h107d9, 'h107e9, 'h10a46, 'h107f9, 'h10809, 'h10a47, 'h103bc, 'h10819, 'h10829, 'h10a48, 'h21f8e, 'h21f8f, 'h21f8d, 'h10839, 'h10849, 'h10a49, 'h10c49, 'h10859, 'h10869, 'h10a4a, 'h10879, 'h10889, 'h10a4b, 'h10899, 'h108a9, 'h10a4c, 'h108b9, 'h103bc, 'h108c9, 'h10a4d, 'h108d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e9, 'h10a4e, 'h10c59, 'h106f9, 'h10709, 'h10a4f, 'h10719, 'h10729, 'h10a50, 'h10739, 'h10749, 'h10a51, 'h10759, 'h10769, 'h10a52, 'h103bc, 'h10779, 'h10789, 'h10a53, 'h21f8e, 'h21f8f, 'h21f8d, 'h10799, 'h10c59, 'h107a9, 'h10a54, 'h107b9, 'h107c9, 'h10a55, 'h107d9, 'h107e9, 'h10a56, 'h107f9, 'h10809, 'h10a57, 'h10819, 'h103bc, 'h10829, 'h10a58, 'h10839, 'h21f8e, 'h21f8f, 'h21f8d, 'h10849, 'h10a59, 'h10c59, 'h10859, 'h10869, 'h10a5a, 'h10879, 'h10889, 'h10a5b, 'h10899, 'h108a9, 'h10a5c, 'h108b9, 'h108c9, 'h10a5d, 'h103bc, 'h108d9, 'h106e9, 'h10a5e, 'h10c69, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f9, 'h10709, 'h10a5f, 'h10719, 'h10729, 'h10a60, 'h10739, 'h10749, 'h10a61, 'h10759, 'h10769, 'h10a62, 'h10779, 'h103bc, 'h10789, 'h10a63, 'h10799, 'h10c69, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a9, 'h10a64, 'h107b9, 'h107c9, 'h10a65, 'h107d9, 'h107e9, 'h10a66, 'h107f9, 'h10809, 'h10a67, 'h10819, 'h10829, 'h10a68, 'h103bc, 'h10839, 'h10849, 'h10a69, 'h10c69, 'h21f8e, 'h21f8f, 'h21f8d, 'h10859, 'h10869, 'h10a6a, 'h10879, 'h10889, 'h10a6b, 'h10899, 'h108a9, 'h10a6c, 'h108b9, 'h108c9, 'h10a6d, 'h108d9, 'h103bc, 'h106e9, 'h10a6e, 'h10c79, 'h106f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10a6f, 'h10719, 'h10729, 'h10a70, 'h10739, 'h10749, 'h10a71, 'h10759, 'h10769, 'h10a72, 'h10779, 'h10789, 'h10a73, 'h103bc, 'h10799, 'h10c79, 'h107a9, 'h10a74, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b9, 'h107c9, 'h10a75, 'h107d9, 'h107e9, 'h10a76, 'h107f9, 'h10809, 'h10a77, 'h10819, 'h10829, 'h10a78, 'h10839, 'h103bc, 'h10849, 'h10a79, 'h10c79, 'h10859, 'h21f8e, 'h21f8f, 'h21f8d, 'h10869, 'h10a7a, 'h10879, 'h10889, 'h10a7b, 'h10899, 'h108a9, 'h10a7c, 'h108b9, 'h108c9, 'h10a7d, 'h108d9, 'h106e9, 'h10a7e, 'h10c89, 'h103bc, 'h106f9, 'h10709, 'h10a7f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10719, 'h10729, 'h10a80, 'h10739, 'h10749, 'h10a81, 'h10759, 'h10769, 'h10a82, 'h10779, 'h10789, 'h10a83, 'h10799, 'h10c89, 'h103bc, 'h107a9, 'h10a84, 'h107b9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c9, 'h10a85, 'h107d9, 'h107e9, 'h10a86, 'h107f9, 'h10809, 'h10a87, 'h10819, 'h10829, 'h10a88, 'h10839, 'h10849, 'h10a89, 'h10c89, 'h103bc, 'h10859, 'h10869, 'h10a8a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10879, 'h10889, 'h10a8b, 'h10899, 'h108a9, 'h10a8c, 'h108b9, 'h108c9, 'h10a8d, 'h108d9, 'h106e9, 'h10a8e, 'h10c99, 'h106f9, 'h103bc, 'h10709, 'h10a8f, 'h10719, 'h21f8e, 'h21f8f, 'h21f8d, 'h10729, 'h10a90, 'h10739, 'h10749, 'h10a91, 'h10759, 'h10769, 'h10a92, 'h10779, 'h10789, 'h10a93, 'h10799, 'h10c99, 'h107a9, 'h10a94, 'h103bc, 'h107b9, 'h107c9, 'h10a95, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d9, 'h107e9, 'h10a96, 'h107f9, 'h10809, 'h10a97, 'h10819, 'h10829, 'h10a98, 'h10839, 'h10849, 'h10a99, 'h10c99, 'h10859, 'h103bc, 'h10869, 'h10a9a, 'h10879, 'h21f8e, 'h21f8f, 'h21f8d, 'h10889, 'h10a9b, 'h10899, 'h108a9, 'h10a9c, 'h108b9, 'h108c9, 'h10a9d, 'h108d9, 'h106e9, 'h10a9e, 'h10ca9, 'h106f9, 'h10709, 'h10a9f, 'h103bc, 'h10719, 'h10729, 'h10aa0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10749, 'h10aa1, 'h10759, 'h10769, 'h10aa2, 'h10779, 'h10789, 'h10aa3, 'h10799, 'h10ca9, 'h107a9, 'h10aa4, 'h107b9, 'h103bc, 'h107c9, 'h10aa5, 'h107d9, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e9, 'h10aa6, 'h107f9, 'h10809, 'h10aa7, 'h10819, 'h10829, 'h10aa8, 'h10839, 'h10849, 'h10aa9, 'h10ca9, 'h10859, 'h10869, 'h10aaa, 'h103bc, 'h10879, 'h10889, 'h10aab, 'h21f8e, 'h21f8f, 'h21f8d, 'h10899, 'h108a9, 'h10aac, 'h108b9, 'h108c9, 'h10aad, 'h108d9, 'h106e9, 'h10aae, 'h10cb9, 'h106f9, 'h10709, 'h10aaf, 'h10719, 'h103bc, 'h10729, 'h10ab0, 'h10739, 'h21f8e, 'h21f8f, 'h21f8d, 'h10749, 'h10ab1, 'h10759, 'h10769, 'h10ab2, 'h10779, 'h10789, 'h10ab3, 'h10799, 'h10cb9, 'h107a9, 'h10ab4, 'h107b9, 'h107c9, 'h10ab5, 'h103bc, 'h107d9, 'h107e9, 'h10ab6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f9, 'h10809, 'h10ab7, 'h10819, 'h10829, 'h10ab8, 'h10839, 'h10849, 'h10ab9, 'h10cb9, 'h10859, 'h10869, 'h10aba, 'h10879, 'h103bc, 'h10889, 'h10abb, 'h10899, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a9, 'h10abc, 'h108b9, 'h108c9, 'h10abd, 'h108d9, 'h106e9, 'h10abe, 'h10cc9, 'h106f9, 'h10709, 'h10abf, 'h10719, 'h10729, 'h10ac0, 'h103bc, 'h10739, 'h10749, 'h10ac1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10759, 'h10769, 'h10ac2, 'h10779, 'h10789, 'h10ac3, 'h10799, 'h10cc9, 'h107a9, 'h10ac4, 'h107b9, 'h107c9, 'h10ac5, 'h107d9, 'h103bc, 'h107e9, 'h10ac6, 'h107f9, 'h21f8e, 'h21f8f, 'h21f8d, 'h10809, 'h10ac7, 'h10819, 'h10829, 'h10ac8, 'h10839};
	int DATA6 [6*SIZE-1:0] = {DATA5, DATA0};
	
endpackage
