

package MATRIX_MULTIPLY_32_PKG_3;
	
	import MATRIX_MULTIPLY_32_PKG_2::DATA2;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h10891, 'h108a1, 'h10adc, 'h108b1, 'h108c1, 'h10add, 'h108d1, 'h106e1, 'h108de, 'h10ae1, 'h106f1, 'h103bc, 'h10701, 'h108df, 'h10711, 'h21f8e, 'h21f8f, 'h21f8d, 'h10721, 'h108e0, 'h10731, 'h10741, 'h108e1, 'h10751, 'h10761, 'h108e2, 'h10771, 'h10781, 'h108e3, 'h10791, 'h10ae1, 'h107a1, 'h108e4, 'h103bc, 'h107b1, 'h107c1, 'h108e5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d1, 'h107e1, 'h108e6, 'h107f1, 'h10801, 'h108e7, 'h10811, 'h10821, 'h108e8, 'h10831, 'h10841, 'h108e9, 'h10ae1, 'h10851, 'h103bc, 'h10861, 'h108ea, 'h10871, 'h21f8e, 'h21f8f, 'h21f8d, 'h10881, 'h108eb, 'h10891, 'h108a1, 'h108ec, 'h108b1, 'h108c1, 'h108ed, 'h108d1, 'h106e1, 'h108ee, 'h10af1, 'h106f1, 'h10701, 'h108ef, 'h103bc, 'h10711, 'h10721, 'h108f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10731, 'h10741, 'h108f1, 'h10751, 'h10761, 'h108f2, 'h10771, 'h10781, 'h108f3, 'h10791, 'h10af1, 'h107a1, 'h108f4, 'h107b1, 'h103bc, 'h107c1, 'h108f5, 'h107d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e1, 'h108f6, 'h107f1, 'h10801, 'h108f7, 'h10811, 'h10821, 'h108f8, 'h10831, 'h10841, 'h108f9, 'h10af1, 'h10851, 'h10861, 'h108fa, 'h103bc, 'h10871, 'h10881, 'h108fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10891, 'h108a1, 'h108fc, 'h108b1, 'h108c1, 'h108fd, 'h108d1, 'h106e1, 'h108fe, 'h10b01, 'h106f1, 'h10701, 'h108ff, 'h10711, 'h103bc, 'h10721, 'h10900, 'h10731, 'h21f8e, 'h21f8f, 'h21f8d, 'h10741, 'h10901, 'h10751, 'h10761, 'h10902, 'h10771, 'h10781, 'h10903, 'h10791, 'h10b01, 'h107a1, 'h10904, 'h107b1, 'h107c1, 'h10905, 'h103bc, 'h107d1, 'h107e1, 'h10906, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f1, 'h10801, 'h10907, 'h10811, 'h10821, 'h10908, 'h10831, 'h10841, 'h10909, 'h10b01, 'h10851, 'h10861, 'h1090a, 'h10871, 'h103bc, 'h10881, 'h1090b, 'h10891, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a1, 'h1090c, 'h108b1, 'h108c1, 'h1090d, 'h108d1, 'h106e1, 'h1090e, 'h10b11, 'h106f1, 'h10701, 'h1090f, 'h10711, 'h10721, 'h10910, 'h103bc, 'h10731, 'h10741, 'h10911, 'h21f8e, 'h21f8f, 'h21f8d, 'h10751, 'h10761, 'h10912, 'h10771, 'h10781, 'h10913, 'h10791, 'h10b11, 'h107a1, 'h10914, 'h107b1, 'h107c1, 'h10915, 'h107d1, 'h103bc, 'h107e1, 'h10916, 'h107f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10801, 'h10917, 'h10811, 'h10821, 'h10918, 'h10831, 'h10841, 'h10919, 'h10b11, 'h10851, 'h10861, 'h1091a, 'h10871, 'h10881, 'h1091b, 'h103bc, 'h10891, 'h108a1, 'h1091c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b1, 'h108c1, 'h1091d, 'h108d1, 'h106e1, 'h1091e, 'h10b21, 'h106f1, 'h10701, 'h1091f, 'h10711, 'h10721, 'h10920, 'h10731, 'h103bc, 'h10741, 'h10921, 'h10751, 'h21f8e, 'h21f8f, 'h21f8d, 'h10761, 'h10922, 'h10771, 'h10781, 'h10923, 'h10791, 'h10b21, 'h107a1, 'h10924, 'h107b1, 'h107c1, 'h10925, 'h107d1, 'h107e1, 'h10926, 'h103bc, 'h107f1, 'h10801, 'h10927, 'h21f8e, 'h21f8f, 'h21f8d, 'h10811, 'h10821, 'h10928, 'h10831, 'h10841, 'h10929, 'h10b21, 'h10851, 'h10861, 'h1092a, 'h10871, 'h10881, 'h1092b, 'h10891, 'h103bc, 'h108a1, 'h1092c, 'h108b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c1, 'h1092d, 'h108d1, 'h106e1, 'h1092e, 'h10b31, 'h106f1, 'h10701, 'h1092f, 'h10711, 'h10721, 'h10930, 'h10731, 'h10741, 'h10931, 'h103bc, 'h10751, 'h10761, 'h10932, 'h21f8e, 'h21f8f, 'h21f8d, 'h10771, 'h10781, 'h10933, 'h10791, 'h10b31, 'h107a1, 'h10934, 'h107b1, 'h107c1, 'h10935, 'h107d1, 'h107e1, 'h10936, 'h107f1, 'h103bc, 'h10801, 'h10937, 'h10811, 'h21f8e, 'h21f8f, 'h21f8d, 'h10821, 'h10938, 'h10831, 'h10841, 'h10939, 'h10b31, 'h10851, 'h10861, 'h1093a, 'h10871, 'h10881, 'h1093b, 'h10891, 'h108a1, 'h1093c, 'h103bc, 'h108b1, 'h108c1, 'h1093d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d1, 'h106e1, 'h1093e, 'h10b41, 'h106f1, 'h10701, 'h1093f, 'h10711, 'h10721, 'h10940, 'h10731, 'h10741, 'h10941, 'h10751, 'h103bc, 'h10761, 'h10942, 'h10771, 'h21f8e, 'h21f8f, 'h21f8d, 'h10781, 'h10943, 'h10791, 'h10b41, 'h107a1, 'h10944, 'h107b1, 'h107c1, 'h10945, 'h107d1, 'h107e1, 'h10946, 'h107f1, 'h10801, 'h10947, 'h103bc, 'h10811, 'h10821, 'h10948, 'h21f8e, 'h21f8f, 'h21f8d, 'h10831, 'h10841, 'h10949, 'h10b41, 'h10851, 'h10861, 'h1094a, 'h10871, 'h10881, 'h1094b, 'h10891, 'h108a1, 'h1094c, 'h108b1, 'h103bc, 'h108c1, 'h1094d, 'h108d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1094e, 'h10b51, 'h106f1, 'h10701, 'h1094f, 'h10711, 'h10721, 'h10950, 'h10731, 'h10741, 'h10951, 'h10751, 'h10761, 'h10952, 'h103bc, 'h10771, 'h10781, 'h10953, 'h21f8e, 'h21f8f, 'h21f8d, 'h10791, 'h10b51, 'h107a1, 'h10954, 'h107b1, 'h107c1, 'h10955, 'h107d1, 'h107e1, 'h10956, 'h107f1, 'h10801, 'h10957, 'h10811, 'h103bc, 'h10821, 'h10958, 'h10831, 'h21f8e, 'h21f8f, 'h21f8d, 'h10841, 'h10959, 'h10b51, 'h10851, 'h10861, 'h1095a, 'h10871, 'h10881, 'h1095b, 'h10891, 'h108a1, 'h1095c, 'h108b1, 'h108c1, 'h1095d, 'h103bc, 'h108d1, 'h106e1, 'h1095e, 'h10b61, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f1, 'h10701, 'h1095f, 'h10711, 'h10721, 'h10960, 'h10731, 'h10741, 'h10961, 'h10751, 'h10761, 'h10962, 'h10771, 'h103bc, 'h10781, 'h10963, 'h10791, 'h10b61, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a1, 'h10964, 'h107b1, 'h107c1, 'h10965, 'h107d1, 'h107e1, 'h10966, 'h107f1, 'h10801, 'h10967, 'h10811, 'h10821, 'h10968, 'h103bc, 'h10831, 'h10841, 'h10969, 'h10b61, 'h21f8e, 'h21f8f, 'h21f8d, 'h10851, 'h10861, 'h1096a, 'h10871, 'h10881, 'h1096b, 'h10891, 'h108a1, 'h1096c, 'h108b1, 'h108c1, 'h1096d, 'h108d1, 'h103bc, 'h106e1, 'h1096e, 'h10b71, 'h106f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10701, 'h1096f, 'h10711, 'h10721, 'h10970, 'h10731, 'h10741, 'h10971, 'h10751, 'h10761, 'h10972, 'h10771, 'h10781, 'h10973, 'h103bc, 'h10791, 'h10b71, 'h107a1, 'h10974, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b1, 'h107c1, 'h10975, 'h107d1, 'h107e1, 'h10976, 'h107f1, 'h10801, 'h10977, 'h10811, 'h10821, 'h10978, 'h10831, 'h103bc, 'h10841, 'h10979, 'h10b71, 'h10851, 'h21f8e, 'h21f8f, 'h21f8d, 'h10861, 'h1097a, 'h10871, 'h10881, 'h1097b, 'h10891, 'h108a1, 'h1097c, 'h108b1, 'h108c1, 'h1097d, 'h108d1, 'h106e1, 'h1097e, 'h10b81, 'h103bc, 'h106f1, 'h10701, 'h1097f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10711, 'h10721, 'h10980, 'h10731, 'h10741, 'h10981, 'h10751, 'h10761, 'h10982, 'h10771, 'h10781, 'h10983, 'h10791, 'h10b81, 'h103bc, 'h107a1, 'h10984, 'h107b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c1, 'h10985, 'h107d1, 'h107e1, 'h10986, 'h107f1, 'h10801, 'h10987, 'h10811, 'h10821, 'h10988, 'h10831, 'h10841, 'h10989, 'h10b81, 'h103bc, 'h10851, 'h10861, 'h1098a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10871, 'h10881, 'h1098b, 'h10891, 'h108a1, 'h1098c, 'h108b1, 'h108c1, 'h1098d, 'h108d1, 'h106e1, 'h1098e, 'h10b91, 'h106f1, 'h103bc, 'h10701, 'h1098f, 'h10711, 'h21f8e, 'h21f8f, 'h21f8d, 'h10721, 'h10990, 'h10731, 'h10741, 'h10991, 'h10751, 'h10761, 'h10992, 'h10771, 'h10781, 'h10993, 'h10791, 'h10b91, 'h107a1, 'h10994, 'h103bc, 'h107b1, 'h107c1, 'h10995, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d1, 'h107e1, 'h10996, 'h107f1, 'h10801, 'h10997, 'h10811, 'h10821, 'h10998, 'h10831, 'h10841, 'h10999, 'h10b91, 'h10851, 'h103bc, 'h10861, 'h1099a, 'h10871, 'h21f8e, 'h21f8f, 'h21f8d, 'h10881, 'h1099b, 'h10891, 'h108a1, 'h1099c, 'h108b1, 'h108c1, 'h1099d, 'h108d1, 'h106e1, 'h1099e, 'h10ba1, 'h106f1, 'h10701, 'h1099f, 'h103bc, 'h10711, 'h10721, 'h109a0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10731, 'h10741, 'h109a1, 'h10751, 'h10761, 'h109a2, 'h10771, 'h10781, 'h109a3, 'h10791, 'h10ba1, 'h107a1, 'h109a4, 'h107b1, 'h103bc, 'h107c1, 'h109a5, 'h107d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e1, 'h109a6, 'h107f1, 'h10801, 'h109a7, 'h10811, 'h10821, 'h109a8, 'h10831, 'h10841, 'h109a9, 'h10ba1, 'h10851, 'h10861, 'h109aa, 'h103bc, 'h10871, 'h10881, 'h109ab, 'h21f8e, 'h21f8f, 'h21f8d, 'h10891, 'h108a1, 'h109ac, 'h108b1, 'h108c1, 'h109ad, 'h108d1, 'h106e1, 'h109ae, 'h10bb1, 'h106f1, 'h10701, 'h109af, 'h10711, 'h103bc, 'h10721, 'h109b0, 'h10731, 'h21f8e, 'h21f8f, 'h21f8d, 'h10741, 'h109b1, 'h10751, 'h10761, 'h109b2, 'h10771, 'h10781, 'h109b3, 'h10791, 'h10bb1, 'h107a1, 'h109b4, 'h107b1, 'h107c1, 'h109b5, 'h103bc, 'h107d1, 'h107e1, 'h109b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f1, 'h10801, 'h109b7, 'h10811, 'h10821, 'h109b8, 'h10831, 'h10841, 'h109b9, 'h10bb1, 'h10851, 'h10861, 'h109ba, 'h10871, 'h103bc, 'h10881, 'h109bb, 'h10891, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a1, 'h109bc, 'h108b1, 'h108c1, 'h109bd, 'h108d1, 'h106e1, 'h109be, 'h10bc1, 'h106f1, 'h10701, 'h109bf, 'h10711, 'h10721, 'h109c0, 'h103bc, 'h10731, 'h10741, 'h109c1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10751, 'h10761, 'h109c2, 'h10771, 'h10781, 'h109c3, 'h10791, 'h10bc1, 'h107a1, 'h109c4, 'h107b1, 'h107c1, 'h109c5, 'h107d1, 'h103bc, 'h107e1, 'h109c6, 'h107f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10801, 'h109c7, 'h10811, 'h10821, 'h109c8, 'h10831, 'h10841, 'h109c9, 'h10bc1, 'h10851, 'h10861, 'h109ca, 'h10871, 'h10881, 'h109cb, 'h103bc, 'h10891, 'h108a1, 'h109cc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b1, 'h108c1, 'h109cd, 'h108d1, 'h106e1, 'h109ce, 'h10bd1, 'h106f1, 'h10701, 'h109cf, 'h10711, 'h10721, 'h109d0, 'h10731, 'h103bc, 'h10741, 'h109d1, 'h10751, 'h21f8e, 'h21f8f, 'h21f8d, 'h10761, 'h109d2, 'h10771, 'h10781, 'h109d3, 'h10791, 'h10bd1, 'h107a1, 'h109d4, 'h107b1, 'h107c1, 'h109d5, 'h107d1, 'h107e1, 'h109d6, 'h103bc, 'h107f1, 'h10801, 'h109d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10811, 'h10821, 'h109d8, 'h10831, 'h10841, 'h109d9, 'h10bd1, 'h10851, 'h10861, 'h109da, 'h10871, 'h10881, 'h109db, 'h10891, 'h103bc, 'h108a1, 'h109dc, 'h108b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c1, 'h109dd, 'h108d1, 'h106e1, 'h109de, 'h10be1, 'h106f1, 'h10701, 'h109df, 'h10711, 'h10721, 'h109e0, 'h10731, 'h10741, 'h109e1, 'h103bc, 'h10751, 'h10761, 'h109e2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10771, 'h10781, 'h109e3, 'h10791, 'h10be1, 'h107a1, 'h109e4, 'h107b1, 'h107c1, 'h109e5, 'h107d1, 'h107e1, 'h109e6, 'h107f1, 'h103bc, 'h10801, 'h109e7, 'h10811, 'h21f8e, 'h21f8f, 'h21f8d, 'h10821, 'h109e8, 'h10831, 'h10841, 'h109e9, 'h10be1, 'h10851, 'h10861, 'h109ea, 'h10871, 'h10881, 'h109eb, 'h10891, 'h108a1, 'h109ec, 'h103bc, 'h108b1, 'h108c1, 'h109ed, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d1, 'h106e1, 'h109ee, 'h10bf1, 'h106f1, 'h10701, 'h109ef, 'h10711, 'h10721, 'h109f0, 'h10731, 'h10741, 'h109f1, 'h10751, 'h103bc, 'h10761, 'h109f2, 'h10771, 'h21f8e, 'h21f8f, 'h21f8d, 'h10781, 'h109f3, 'h10791, 'h10bf1, 'h107a1, 'h109f4, 'h107b1, 'h107c1, 'h109f5, 'h107d1, 'h107e1, 'h109f6, 'h107f1, 'h10801, 'h109f7, 'h103bc, 'h10811, 'h10821, 'h109f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10831, 'h10841, 'h109f9, 'h10bf1, 'h10851, 'h10861, 'h109fa, 'h10871, 'h10881, 'h109fb, 'h10891, 'h108a1, 'h109fc, 'h108b1, 'h103bc, 'h108c1, 'h109fd, 'h108d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h109fe, 'h10c01, 'h106f1, 'h10701, 'h109ff, 'h10711, 'h10721, 'h10a00, 'h10731, 'h10741, 'h10a01, 'h10751, 'h10761, 'h10a02, 'h103bc, 'h10771, 'h10781, 'h10a03, 'h21f8e, 'h21f8f, 'h21f8d, 'h10791, 'h10c01, 'h107a1, 'h10a04, 'h107b1, 'h107c1, 'h10a05, 'h107d1, 'h107e1, 'h10a06, 'h107f1, 'h10801, 'h10a07, 'h10811, 'h103bc, 'h10821, 'h10a08, 'h10831, 'h21f8e, 'h21f8f, 'h21f8d, 'h10841, 'h10a09, 'h10c01, 'h10851, 'h10861, 'h10a0a, 'h10871, 'h10881, 'h10a0b, 'h10891, 'h108a1, 'h10a0c, 'h108b1, 'h108c1, 'h10a0d, 'h103bc, 'h108d1, 'h106e1, 'h10a0e, 'h10c11, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f1, 'h10701, 'h10a0f, 'h10711, 'h10721, 'h10a10, 'h10731, 'h10741, 'h10a11, 'h10751, 'h10761, 'h10a12, 'h10771, 'h103bc, 'h10781, 'h10a13, 'h10791, 'h10c11, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a1, 'h10a14, 'h107b1, 'h107c1, 'h10a15, 'h107d1, 'h107e1, 'h10a16, 'h107f1, 'h10801, 'h10a17, 'h10811, 'h10821, 'h10a18, 'h103bc, 'h10831, 'h10841, 'h10a19, 'h10c11, 'h21f8e, 'h21f8f, 'h21f8d, 'h10851, 'h10861, 'h10a1a, 'h10871, 'h10881, 'h10a1b, 'h10891, 'h108a1, 'h10a1c, 'h108b1, 'h108c1, 'h10a1d, 'h108d1, 'h103bc, 'h106e1, 'h10a1e, 'h10c21, 'h106f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10701, 'h10a1f, 'h10711, 'h10721, 'h10a20, 'h10731, 'h10741, 'h10a21, 'h10751, 'h10761, 'h10a22, 'h10771, 'h10781, 'h10a23, 'h103bc, 'h10791, 'h10c21, 'h107a1, 'h10a24, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b1, 'h107c1, 'h10a25, 'h107d1, 'h107e1, 'h10a26, 'h107f1, 'h10801, 'h10a27, 'h10811, 'h10821, 'h10a28, 'h10831, 'h103bc, 'h10841, 'h10a29, 'h10c21, 'h10851, 'h21f8e, 'h21f8f, 'h21f8d, 'h10861, 'h10a2a, 'h10871, 'h10881, 'h10a2b, 'h10891, 'h108a1, 'h10a2c, 'h108b1, 'h108c1, 'h10a2d, 'h108d1, 'h106e1, 'h10a2e, 'h10c31, 'h103bc, 'h106f1, 'h10701, 'h10a2f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10711, 'h10721, 'h10a30, 'h10731, 'h10741, 'h10a31, 'h10751, 'h10761, 'h10a32, 'h10771, 'h10781, 'h10a33, 'h10791, 'h10c31, 'h103bc, 'h107a1, 'h10a34, 'h107b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c1, 'h10a35, 'h107d1, 'h107e1, 'h10a36, 'h107f1, 'h10801, 'h10a37, 'h10811, 'h10821, 'h10a38, 'h10831, 'h10841, 'h10a39, 'h10c31, 'h103bc, 'h10851, 'h10861, 'h10a3a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10871, 'h10881, 'h10a3b, 'h10891, 'h108a1, 'h10a3c, 'h108b1, 'h108c1, 'h10a3d, 'h108d1, 'h106e1, 'h10a3e, 'h10c41, 'h106f1, 'h103bc, 'h10701, 'h10a3f, 'h10711, 'h21f8e, 'h21f8f, 'h21f8d, 'h10721, 'h10a40, 'h10731, 'h10741, 'h10a41, 'h10751, 'h10761, 'h10a42, 'h10771, 'h10781, 'h10a43, 'h10791, 'h10c41, 'h107a1, 'h10a44, 'h103bc, 'h107b1, 'h107c1, 'h10a45, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d1, 'h107e1, 'h10a46, 'h107f1, 'h10801, 'h10a47, 'h10811, 'h10821, 'h10a48, 'h10831, 'h10841, 'h10a49, 'h10c41, 'h10851, 'h103bc, 'h10861, 'h10a4a, 'h10871, 'h21f8e, 'h21f8f, 'h21f8d, 'h10881, 'h10a4b, 'h10891, 'h108a1, 'h10a4c, 'h108b1, 'h108c1, 'h10a4d, 'h108d1, 'h106e1, 'h10a4e, 'h10c51, 'h106f1, 'h10701, 'h10a4f, 'h103bc, 'h10711, 'h10721, 'h10a50, 'h21f8e, 'h21f8f, 'h21f8d, 'h10731, 'h10741, 'h10a51, 'h10751, 'h10761, 'h10a52, 'h10771, 'h10781, 'h10a53, 'h10791, 'h10c51, 'h107a1, 'h10a54, 'h107b1, 'h103bc, 'h107c1, 'h10a55, 'h107d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e1, 'h10a56, 'h107f1, 'h10801, 'h10a57, 'h10811, 'h10821, 'h10a58, 'h10831, 'h10841, 'h10a59, 'h10c51, 'h10851, 'h10861, 'h10a5a, 'h103bc, 'h10871, 'h10881, 'h10a5b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10891, 'h108a1, 'h10a5c, 'h108b1, 'h108c1, 'h10a5d, 'h108d1, 'h106e1, 'h10a5e, 'h10c61, 'h106f1, 'h10701, 'h10a5f, 'h10711, 'h103bc, 'h10721, 'h10a60, 'h10731, 'h21f8e, 'h21f8f, 'h21f8d, 'h10741, 'h10a61, 'h10751, 'h10761, 'h10a62, 'h10771, 'h10781, 'h10a63, 'h10791, 'h10c61, 'h107a1, 'h10a64, 'h107b1, 'h107c1, 'h10a65, 'h103bc, 'h107d1, 'h107e1, 'h10a66, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f1, 'h10801, 'h10a67, 'h10811, 'h10821, 'h10a68, 'h10831, 'h10841, 'h10a69, 'h10c61, 'h10851, 'h10861, 'h10a6a, 'h10871, 'h103bc, 'h10881, 'h10a6b, 'h10891, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a1, 'h10a6c, 'h108b1, 'h108c1, 'h10a6d, 'h108d1, 'h106e1, 'h10a6e, 'h10c71, 'h106f1, 'h10701, 'h10a6f, 'h10711, 'h10721, 'h10a70, 'h103bc, 'h10731, 'h10741, 'h10a71, 'h21f8e, 'h21f8f, 'h21f8d, 'h10751, 'h10761, 'h10a72, 'h10771, 'h10781, 'h10a73, 'h10791, 'h10c71, 'h107a1, 'h10a74, 'h107b1, 'h107c1, 'h10a75, 'h107d1, 'h103bc, 'h107e1, 'h10a76, 'h107f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10801, 'h10a77, 'h10811, 'h10821, 'h10a78, 'h10831, 'h10841, 'h10a79, 'h10c71, 'h10851, 'h10861, 'h10a7a, 'h10871, 'h10881, 'h10a7b, 'h103bc, 'h10891, 'h108a1, 'h10a7c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b1, 'h108c1, 'h10a7d, 'h108d1, 'h106e1, 'h10a7e, 'h10c81, 'h106f1, 'h10701, 'h10a7f, 'h10711, 'h10721, 'h10a80, 'h10731, 'h103bc, 'h10741, 'h10a81, 'h10751, 'h21f8e, 'h21f8f, 'h21f8d, 'h10761, 'h10a82, 'h10771, 'h10781, 'h10a83, 'h10791, 'h10c81, 'h107a1, 'h10a84, 'h107b1, 'h107c1, 'h10a85, 'h107d1, 'h107e1, 'h10a86, 'h103bc, 'h107f1, 'h10801, 'h10a87, 'h21f8e, 'h21f8f, 'h21f8d, 'h10811, 'h10821, 'h10a88, 'h10831, 'h10841, 'h10a89, 'h10c81, 'h10851, 'h10861, 'h10a8a, 'h10871, 'h10881, 'h10a8b, 'h10891, 'h103bc, 'h108a1, 'h10a8c, 'h108b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c1, 'h10a8d, 'h108d1, 'h106e1, 'h10a8e, 'h10c91, 'h106f1, 'h10701, 'h10a8f, 'h10711, 'h10721, 'h10a90, 'h10731, 'h10741, 'h10a91, 'h103bc, 'h10751, 'h10761, 'h10a92, 'h21f8e, 'h21f8f, 'h21f8d, 'h10771, 'h10781, 'h10a93, 'h10791, 'h10c91, 'h107a1, 'h10a94, 'h107b1, 'h107c1, 'h10a95, 'h107d1, 'h107e1, 'h10a96, 'h107f1, 'h103bc, 'h10801, 'h10a97, 'h10811, 'h21f8e, 'h21f8f, 'h21f8d, 'h10821, 'h10a98, 'h10831, 'h10841, 'h10a99, 'h10c91, 'h10851, 'h10861, 'h10a9a, 'h10871, 'h10881, 'h10a9b, 'h10891, 'h108a1, 'h10a9c, 'h103bc, 'h108b1, 'h108c1, 'h10a9d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d1, 'h106e1, 'h10a9e, 'h10ca1, 'h106f1, 'h10701, 'h10a9f, 'h10711, 'h10721, 'h10aa0, 'h10731, 'h10741, 'h10aa1, 'h10751, 'h103bc, 'h10761, 'h10aa2, 'h10771, 'h21f8e, 'h21f8f, 'h21f8d, 'h10781, 'h10aa3, 'h10791, 'h10ca1, 'h107a1, 'h10aa4, 'h107b1, 'h107c1, 'h10aa5, 'h107d1, 'h107e1, 'h10aa6, 'h107f1, 'h10801, 'h10aa7, 'h103bc, 'h10811, 'h10821, 'h10aa8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10831, 'h10841, 'h10aa9, 'h10ca1, 'h10851, 'h10861, 'h10aaa, 'h10871, 'h10881, 'h10aab, 'h10891, 'h108a1, 'h10aac, 'h108b1, 'h103bc, 'h108c1, 'h10aad, 'h108d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h10aae, 'h10cb1, 'h106f1, 'h10701, 'h10aaf, 'h10711, 'h10721, 'h10ab0, 'h10731, 'h10741, 'h10ab1, 'h10751, 'h10761, 'h10ab2, 'h103bc, 'h10771, 'h10781, 'h10ab3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10791, 'h10cb1, 'h107a1, 'h10ab4, 'h107b1, 'h107c1, 'h10ab5, 'h107d1, 'h107e1, 'h10ab6, 'h107f1, 'h10801, 'h10ab7, 'h10811, 'h103bc, 'h10821, 'h10ab8, 'h10831, 'h21f8e, 'h21f8f, 'h21f8d, 'h10841, 'h10ab9, 'h10cb1, 'h10851, 'h10861, 'h10aba, 'h10871, 'h10881, 'h10abb, 'h10891, 'h108a1, 'h10abc, 'h108b1, 'h108c1, 'h10abd, 'h103bc, 'h108d1, 'h106e1, 'h10abe, 'h10cc1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f1, 'h10701, 'h10abf, 'h10711, 'h10721, 'h10ac0, 'h10731, 'h10741, 'h10ac1, 'h10751, 'h10761, 'h10ac2, 'h10771, 'h103bc, 'h10781, 'h10ac3, 'h10791, 'h10cc1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a1, 'h10ac4, 'h107b1, 'h107c1, 'h10ac5, 'h107d1, 'h107e1, 'h10ac6, 'h107f1, 'h10801, 'h10ac7, 'h10811, 'h10821, 'h10ac8, 'h103bc, 'h10831, 'h10841, 'h10ac9, 'h10cc1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10851, 'h10861, 'h10aca, 'h10871, 'h10881, 'h10acb, 'h10891, 'h108a1, 'h10acc, 'h108b1, 'h108c1, 'h10acd, 'h108d1, 'h103bc, 'h106e1, 'h10ace, 'h10cd1, 'h106f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10701, 'h10acf, 'h10711, 'h10721, 'h10ad0, 'h10731, 'h10741, 'h10ad1, 'h10751, 'h10761, 'h10ad2, 'h10771, 'h10781, 'h10ad3, 'h103bc, 'h10791, 'h10cd1, 'h107a1, 'h10ad4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b1, 'h107c1, 'h10ad5, 'h107d1, 'h107e1, 'h10ad6, 'h107f1, 'h10801, 'h10ad7, 'h10811, 'h10821, 'h10ad8, 'h10831, 'h103bc, 'h10841, 'h10ad9, 'h10cd1, 'h10851, 'h21f8e, 'h21f8f, 'h21f8d, 'h10861, 'h10ada, 'h10871, 'h10881, 'h10adb, 'h10891, 'h108a1, 'h10adc, 'h108b1, 'h108c1, 'h10add, 'h108d1, 'h106e2, 'h108de, 'h10ae2, 'h103bc, 'h106f2, 'h10702, 'h108df, 'h21f8e, 'h21f8f, 'h21f8d, 'h10712, 'h10722, 'h108e0, 'h10732, 'h10742, 'h108e1, 'h10752, 'h10762, 'h108e2, 'h10772, 'h10782, 'h108e3, 'h10792, 'h10ae2, 'h103bc, 'h107a2, 'h108e4, 'h107b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c2, 'h108e5, 'h107d2, 'h107e2, 'h108e6, 'h107f2, 'h10802, 'h108e7, 'h10812, 'h10822, 'h108e8, 'h10832, 'h10842, 'h108e9, 'h10ae2, 'h103bc, 'h10852, 'h10862, 'h108ea, 'h21f8e, 'h21f8f, 'h21f8d, 'h10872, 'h10882, 'h108eb, 'h10892, 'h108a2, 'h108ec, 'h108b2, 'h108c2, 'h108ed, 'h108d2, 'h106e2, 'h108ee, 'h10af2, 'h106f2, 'h103bc, 'h10702, 'h108ef, 'h10712, 'h21f8e, 'h21f8f, 'h21f8d, 'h10722, 'h108f0, 'h10732, 'h10742, 'h108f1, 'h10752, 'h10762, 'h108f2, 'h10772, 'h10782, 'h108f3, 'h10792, 'h10af2, 'h107a2, 'h108f4, 'h103bc, 'h107b2, 'h107c2, 'h108f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d2, 'h107e2, 'h108f6, 'h107f2, 'h10802, 'h108f7, 'h10812, 'h10822, 'h108f8, 'h10832, 'h10842, 'h108f9, 'h10af2, 'h10852, 'h103bc, 'h10862, 'h108fa, 'h10872, 'h21f8e, 'h21f8f, 'h21f8d, 'h10882, 'h108fb, 'h10892, 'h108a2, 'h108fc, 'h108b2, 'h108c2, 'h108fd, 'h108d2, 'h106e2, 'h108fe, 'h10b02, 'h106f2, 'h10702, 'h108ff, 'h103bc, 'h10712, 'h10722, 'h10900, 'h21f8e, 'h21f8f, 'h21f8d, 'h10732, 'h10742, 'h10901, 'h10752, 'h10762, 'h10902, 'h10772, 'h10782, 'h10903, 'h10792, 'h10b02, 'h107a2, 'h10904, 'h107b2, 'h103bc, 'h107c2, 'h10905, 'h107d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e2, 'h10906, 'h107f2, 'h10802, 'h10907, 'h10812, 'h10822, 'h10908, 'h10832, 'h10842, 'h10909, 'h10b02, 'h10852, 'h10862, 'h1090a, 'h103bc, 'h10872, 'h10882, 'h1090b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10892, 'h108a2, 'h1090c, 'h108b2, 'h108c2, 'h1090d, 'h108d2, 'h106e2, 'h1090e, 'h10b12, 'h106f2, 'h10702, 'h1090f, 'h10712, 'h103bc, 'h10722, 'h10910, 'h10732, 'h21f8e, 'h21f8f, 'h21f8d, 'h10742, 'h10911, 'h10752, 'h10762, 'h10912, 'h10772, 'h10782, 'h10913, 'h10792, 'h10b12, 'h107a2, 'h10914, 'h107b2, 'h107c2, 'h10915, 'h103bc, 'h107d2, 'h107e2, 'h10916, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f2, 'h10802, 'h10917, 'h10812, 'h10822, 'h10918, 'h10832, 'h10842, 'h10919, 'h10b12, 'h10852, 'h10862, 'h1091a, 'h10872, 'h103bc, 'h10882, 'h1091b, 'h10892, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a2, 'h1091c, 'h108b2, 'h108c2, 'h1091d, 'h108d2, 'h106e2, 'h1091e, 'h10b22, 'h106f2, 'h10702, 'h1091f, 'h10712, 'h10722, 'h10920, 'h103bc, 'h10732, 'h10742, 'h10921, 'h21f8e, 'h21f8f, 'h21f8d, 'h10752, 'h10762, 'h10922, 'h10772, 'h10782, 'h10923, 'h10792, 'h10b22, 'h107a2, 'h10924, 'h107b2, 'h107c2, 'h10925, 'h107d2, 'h103bc, 'h107e2, 'h10926, 'h107f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10802, 'h10927, 'h10812, 'h10822, 'h10928, 'h10832, 'h10842, 'h10929, 'h10b22, 'h10852, 'h10862, 'h1092a, 'h10872, 'h10882, 'h1092b, 'h103bc, 'h10892, 'h108a2, 'h1092c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b2, 'h108c2, 'h1092d, 'h108d2, 'h106e2, 'h1092e, 'h10b32, 'h106f2, 'h10702, 'h1092f, 'h10712, 'h10722, 'h10930, 'h10732, 'h103bc, 'h10742, 'h10931, 'h10752, 'h21f8e, 'h21f8f, 'h21f8d, 'h10762, 'h10932, 'h10772, 'h10782, 'h10933, 'h10792, 'h10b32, 'h107a2, 'h10934, 'h107b2, 'h107c2, 'h10935, 'h107d2, 'h107e2, 'h10936, 'h103bc, 'h107f2, 'h10802, 'h10937, 'h21f8e, 'h21f8f, 'h21f8d, 'h10812, 'h10822, 'h10938, 'h10832, 'h10842, 'h10939, 'h10b32, 'h10852, 'h10862, 'h1093a, 'h10872, 'h10882, 'h1093b, 'h10892, 'h103bc, 'h108a2, 'h1093c, 'h108b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c2, 'h1093d, 'h108d2, 'h106e2, 'h1093e, 'h10b42, 'h106f2, 'h10702, 'h1093f, 'h10712, 'h10722, 'h10940, 'h10732, 'h10742, 'h10941, 'h103bc, 'h10752, 'h10762, 'h10942, 'h21f8e, 'h21f8f, 'h21f8d, 'h10772, 'h10782, 'h10943, 'h10792, 'h10b42, 'h107a2, 'h10944, 'h107b2, 'h107c2, 'h10945, 'h107d2, 'h107e2, 'h10946, 'h107f2, 'h103bc, 'h10802, 'h10947, 'h10812, 'h21f8e, 'h21f8f, 'h21f8d, 'h10822, 'h10948, 'h10832, 'h10842, 'h10949, 'h10b42, 'h10852, 'h10862, 'h1094a, 'h10872, 'h10882, 'h1094b, 'h10892, 'h108a2, 'h1094c, 'h103bc, 'h108b2, 'h108c2, 'h1094d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d2, 'h106e2, 'h1094e, 'h10b52, 'h106f2, 'h10702, 'h1094f, 'h10712, 'h10722, 'h10950, 'h10732, 'h10742, 'h10951, 'h10752, 'h103bc, 'h10762, 'h10952, 'h10772, 'h21f8e, 'h21f8f, 'h21f8d, 'h10782, 'h10953, 'h10792, 'h10b52, 'h107a2, 'h10954, 'h107b2, 'h107c2, 'h10955, 'h107d2, 'h107e2, 'h10956, 'h107f2, 'h10802, 'h10957, 'h103bc, 'h10812, 'h10822, 'h10958, 'h21f8e, 'h21f8f, 'h21f8d, 'h10832, 'h10842, 'h10959, 'h10b52, 'h10852, 'h10862, 'h1095a, 'h10872, 'h10882, 'h1095b, 'h10892, 'h108a2, 'h1095c, 'h108b2, 'h103bc, 'h108c2, 'h1095d, 'h108d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1095e, 'h10b62, 'h106f2, 'h10702, 'h1095f, 'h10712, 'h10722, 'h10960, 'h10732, 'h10742, 'h10961, 'h10752, 'h10762, 'h10962, 'h103bc, 'h10772, 'h10782, 'h10963, 'h21f8e, 'h21f8f, 'h21f8d, 'h10792, 'h10b62, 'h107a2, 'h10964, 'h107b2, 'h107c2, 'h10965, 'h107d2, 'h107e2, 'h10966, 'h107f2, 'h10802, 'h10967, 'h10812, 'h103bc, 'h10822, 'h10968, 'h10832, 'h21f8e, 'h21f8f, 'h21f8d, 'h10842, 'h10969, 'h10b62, 'h10852, 'h10862, 'h1096a, 'h10872, 'h10882, 'h1096b, 'h10892, 'h108a2, 'h1096c, 'h108b2, 'h108c2, 'h1096d, 'h103bc, 'h108d2, 'h106e2, 'h1096e, 'h10b72, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f2, 'h10702, 'h1096f, 'h10712, 'h10722, 'h10970, 'h10732, 'h10742, 'h10971, 'h10752, 'h10762, 'h10972, 'h10772, 'h103bc, 'h10782, 'h10973, 'h10792, 'h10b72, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a2, 'h10974, 'h107b2, 'h107c2, 'h10975, 'h107d2, 'h107e2, 'h10976, 'h107f2, 'h10802, 'h10977, 'h10812, 'h10822, 'h10978, 'h103bc, 'h10832, 'h10842, 'h10979, 'h10b72, 'h21f8e, 'h21f8f, 'h21f8d, 'h10852, 'h10862, 'h1097a, 'h10872, 'h10882, 'h1097b, 'h10892, 'h108a2, 'h1097c, 'h108b2, 'h108c2, 'h1097d, 'h108d2, 'h103bc, 'h106e2, 'h1097e, 'h10b82, 'h106f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10702, 'h1097f, 'h10712, 'h10722, 'h10980, 'h10732, 'h10742, 'h10981, 'h10752, 'h10762, 'h10982, 'h10772, 'h10782, 'h10983, 'h103bc, 'h10792, 'h10b82, 'h107a2, 'h10984, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b2, 'h107c2, 'h10985, 'h107d2, 'h107e2, 'h10986, 'h107f2, 'h10802, 'h10987, 'h10812, 'h10822, 'h10988, 'h10832, 'h103bc, 'h10842, 'h10989, 'h10b82, 'h10852, 'h21f8e, 'h21f8f, 'h21f8d, 'h10862, 'h1098a, 'h10872, 'h10882, 'h1098b, 'h10892, 'h108a2, 'h1098c, 'h108b2, 'h108c2, 'h1098d, 'h108d2, 'h106e2, 'h1098e, 'h10b92, 'h103bc, 'h106f2, 'h10702, 'h1098f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10712, 'h10722, 'h10990, 'h10732, 'h10742, 'h10991, 'h10752, 'h10762, 'h10992, 'h10772, 'h10782, 'h10993, 'h10792, 'h10b92, 'h103bc, 'h107a2, 'h10994, 'h107b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c2, 'h10995, 'h107d2, 'h107e2, 'h10996, 'h107f2, 'h10802, 'h10997, 'h10812, 'h10822, 'h10998, 'h10832, 'h10842, 'h10999, 'h10b92, 'h103bc, 'h10852, 'h10862, 'h1099a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10872, 'h10882, 'h1099b, 'h10892, 'h108a2, 'h1099c, 'h108b2, 'h108c2, 'h1099d, 'h108d2, 'h106e2, 'h1099e, 'h10ba2, 'h106f2, 'h103bc, 'h10702, 'h1099f, 'h10712, 'h21f8e, 'h21f8f, 'h21f8d, 'h10722, 'h109a0, 'h10732, 'h10742, 'h109a1, 'h10752, 'h10762, 'h109a2, 'h10772, 'h10782, 'h109a3, 'h10792, 'h10ba2, 'h107a2, 'h109a4, 'h103bc, 'h107b2, 'h107c2, 'h109a5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d2, 'h107e2, 'h109a6, 'h107f2, 'h10802, 'h109a7, 'h10812, 'h10822, 'h109a8, 'h10832, 'h10842, 'h109a9, 'h10ba2, 'h10852, 'h103bc, 'h10862, 'h109aa, 'h10872, 'h21f8e, 'h21f8f, 'h21f8d, 'h10882, 'h109ab, 'h10892, 'h108a2, 'h109ac, 'h108b2, 'h108c2, 'h109ad, 'h108d2, 'h106e2, 'h109ae, 'h10bb2, 'h106f2, 'h10702, 'h109af, 'h103bc, 'h10712, 'h10722, 'h109b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10732, 'h10742, 'h109b1, 'h10752, 'h10762, 'h109b2, 'h10772, 'h10782, 'h109b3, 'h10792, 'h10bb2, 'h107a2, 'h109b4, 'h107b2, 'h103bc, 'h107c2, 'h109b5, 'h107d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e2, 'h109b6, 'h107f2, 'h10802, 'h109b7, 'h10812, 'h10822, 'h109b8, 'h10832, 'h10842, 'h109b9, 'h10bb2, 'h10852, 'h10862, 'h109ba, 'h103bc, 'h10872, 'h10882, 'h109bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10892, 'h108a2, 'h109bc, 'h108b2, 'h108c2, 'h109bd, 'h108d2, 'h106e2, 'h109be, 'h10bc2, 'h106f2, 'h10702, 'h109bf, 'h10712, 'h103bc, 'h10722, 'h109c0, 'h10732, 'h21f8e, 'h21f8f, 'h21f8d, 'h10742, 'h109c1, 'h10752, 'h10762, 'h109c2, 'h10772, 'h10782, 'h109c3, 'h10792, 'h10bc2, 'h107a2, 'h109c4, 'h107b2, 'h107c2, 'h109c5, 'h103bc, 'h107d2, 'h107e2, 'h109c6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f2, 'h10802, 'h109c7, 'h10812, 'h10822, 'h109c8, 'h10832, 'h10842, 'h109c9, 'h10bc2, 'h10852, 'h10862, 'h109ca, 'h10872, 'h103bc, 'h10882, 'h109cb, 'h10892, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a2, 'h109cc, 'h108b2, 'h108c2, 'h109cd, 'h108d2, 'h106e2, 'h109ce, 'h10bd2, 'h106f2, 'h10702, 'h109cf, 'h10712, 'h10722, 'h109d0, 'h103bc, 'h10732, 'h10742, 'h109d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10752, 'h10762, 'h109d2, 'h10772, 'h10782, 'h109d3, 'h10792, 'h10bd2, 'h107a2, 'h109d4, 'h107b2, 'h107c2, 'h109d5, 'h107d2, 'h103bc, 'h107e2, 'h109d6, 'h107f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10802, 'h109d7, 'h10812, 'h10822, 'h109d8, 'h10832, 'h10842, 'h109d9, 'h10bd2, 'h10852, 'h10862, 'h109da, 'h10872, 'h10882, 'h109db, 'h103bc, 'h10892, 'h108a2, 'h109dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b2, 'h108c2, 'h109dd, 'h108d2, 'h106e2, 'h109de, 'h10be2, 'h106f2, 'h10702, 'h109df, 'h10712, 'h10722, 'h109e0, 'h10732, 'h103bc, 'h10742, 'h109e1, 'h10752, 'h21f8e, 'h21f8f, 'h21f8d, 'h10762, 'h109e2, 'h10772, 'h10782, 'h109e3, 'h10792, 'h10be2, 'h107a2, 'h109e4, 'h107b2, 'h107c2, 'h109e5, 'h107d2, 'h107e2, 'h109e6, 'h103bc, 'h107f2, 'h10802, 'h109e7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10812, 'h10822, 'h109e8, 'h10832, 'h10842, 'h109e9, 'h10be2, 'h10852, 'h10862, 'h109ea, 'h10872, 'h10882, 'h109eb, 'h10892, 'h103bc, 'h108a2, 'h109ec, 'h108b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c2, 'h109ed, 'h108d2, 'h106e2, 'h109ee, 'h10bf2, 'h106f2, 'h10702, 'h109ef, 'h10712, 'h10722, 'h109f0, 'h10732, 'h10742, 'h109f1, 'h103bc, 'h10752, 'h10762, 'h109f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10772, 'h10782, 'h109f3, 'h10792, 'h10bf2, 'h107a2, 'h109f4, 'h107b2, 'h107c2, 'h109f5, 'h107d2, 'h107e2, 'h109f6, 'h107f2, 'h103bc, 'h10802, 'h109f7, 'h10812, 'h21f8e, 'h21f8f, 'h21f8d, 'h10822, 'h109f8, 'h10832, 'h10842, 'h109f9, 'h10bf2, 'h10852, 'h10862, 'h109fa, 'h10872, 'h10882, 'h109fb, 'h10892, 'h108a2, 'h109fc, 'h103bc, 'h108b2, 'h108c2, 'h109fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d2, 'h106e2, 'h109fe, 'h10c02, 'h106f2, 'h10702, 'h109ff, 'h10712, 'h10722, 'h10a00, 'h10732, 'h10742, 'h10a01, 'h10752, 'h103bc, 'h10762, 'h10a02, 'h10772, 'h21f8e, 'h21f8f, 'h21f8d, 'h10782, 'h10a03, 'h10792, 'h10c02, 'h107a2, 'h10a04, 'h107b2, 'h107c2, 'h10a05, 'h107d2, 'h107e2, 'h10a06, 'h107f2, 'h10802, 'h10a07, 'h103bc, 'h10812, 'h10822, 'h10a08, 'h21f8e, 'h21f8f, 'h21f8d, 'h10832, 'h10842, 'h10a09, 'h10c02, 'h10852, 'h10862, 'h10a0a, 'h10872, 'h10882, 'h10a0b, 'h10892, 'h108a2, 'h10a0c, 'h108b2, 'h103bc, 'h108c2, 'h10a0d, 'h108d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h10a0e, 'h10c12, 'h106f2, 'h10702, 'h10a0f, 'h10712, 'h10722, 'h10a10, 'h10732, 'h10742, 'h10a11, 'h10752, 'h10762, 'h10a12, 'h103bc, 'h10772, 'h10782, 'h10a13, 'h21f8e, 'h21f8f, 'h21f8d, 'h10792, 'h10c12, 'h107a2, 'h10a14, 'h107b2, 'h107c2, 'h10a15, 'h107d2, 'h107e2, 'h10a16, 'h107f2, 'h10802, 'h10a17, 'h10812, 'h103bc, 'h10822, 'h10a18, 'h10832, 'h21f8e, 'h21f8f, 'h21f8d, 'h10842, 'h10a19, 'h10c12, 'h10852, 'h10862, 'h10a1a, 'h10872, 'h10882, 'h10a1b, 'h10892, 'h108a2, 'h10a1c, 'h108b2, 'h108c2, 'h10a1d, 'h103bc, 'h108d2, 'h106e2, 'h10a1e, 'h10c22, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f2, 'h10702, 'h10a1f, 'h10712, 'h10722, 'h10a20, 'h10732, 'h10742, 'h10a21, 'h10752, 'h10762, 'h10a22, 'h10772, 'h103bc, 'h10782, 'h10a23, 'h10792, 'h10c22, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a2, 'h10a24, 'h107b2, 'h107c2, 'h10a25, 'h107d2, 'h107e2, 'h10a26, 'h107f2, 'h10802, 'h10a27, 'h10812, 'h10822, 'h10a28, 'h103bc, 'h10832, 'h10842, 'h10a29, 'h10c22, 'h21f8e, 'h21f8f, 'h21f8d, 'h10852, 'h10862, 'h10a2a, 'h10872, 'h10882, 'h10a2b, 'h10892, 'h108a2, 'h10a2c, 'h108b2, 'h108c2, 'h10a2d, 'h108d2, 'h103bc, 'h106e2, 'h10a2e, 'h10c32, 'h106f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10702, 'h10a2f, 'h10712, 'h10722, 'h10a30, 'h10732, 'h10742, 'h10a31, 'h10752, 'h10762, 'h10a32, 'h10772, 'h10782, 'h10a33, 'h103bc, 'h10792, 'h10c32, 'h107a2, 'h10a34, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b2, 'h107c2, 'h10a35, 'h107d2, 'h107e2, 'h10a36, 'h107f2, 'h10802, 'h10a37, 'h10812, 'h10822, 'h10a38, 'h10832, 'h103bc, 'h10842, 'h10a39, 'h10c32, 'h10852, 'h21f8e, 'h21f8f, 'h21f8d, 'h10862, 'h10a3a, 'h10872, 'h10882, 'h10a3b, 'h10892, 'h108a2, 'h10a3c, 'h108b2, 'h108c2, 'h10a3d, 'h108d2, 'h106e2, 'h10a3e, 'h10c42, 'h103bc, 'h106f2, 'h10702, 'h10a3f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10712, 'h10722, 'h10a40, 'h10732, 'h10742, 'h10a41, 'h10752, 'h10762, 'h10a42, 'h10772, 'h10782, 'h10a43, 'h10792, 'h10c42, 'h103bc, 'h107a2, 'h10a44, 'h107b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c2, 'h10a45, 'h107d2, 'h107e2, 'h10a46, 'h107f2, 'h10802, 'h10a47, 'h10812, 'h10822, 'h10a48, 'h10832, 'h10842, 'h10a49, 'h10c42, 'h103bc, 'h10852, 'h10862, 'h10a4a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10872, 'h10882, 'h10a4b, 'h10892, 'h108a2, 'h10a4c, 'h108b2, 'h108c2, 'h10a4d, 'h108d2, 'h106e2, 'h10a4e, 'h10c52, 'h106f2, 'h103bc, 'h10702, 'h10a4f, 'h10712, 'h21f8e, 'h21f8f, 'h21f8d, 'h10722, 'h10a50, 'h10732, 'h10742, 'h10a51, 'h10752, 'h10762, 'h10a52, 'h10772, 'h10782, 'h10a53, 'h10792, 'h10c52, 'h107a2, 'h10a54, 'h103bc, 'h107b2, 'h107c2, 'h10a55, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d2, 'h107e2, 'h10a56, 'h107f2, 'h10802, 'h10a57, 'h10812, 'h10822, 'h10a58, 'h10832, 'h10842, 'h10a59, 'h10c52, 'h10852, 'h103bc, 'h10862, 'h10a5a, 'h10872, 'h21f8e, 'h21f8f, 'h21f8d, 'h10882, 'h10a5b, 'h10892, 'h108a2, 'h10a5c, 'h108b2, 'h108c2, 'h10a5d, 'h108d2, 'h106e2, 'h10a5e, 'h10c62, 'h106f2, 'h10702, 'h10a5f, 'h103bc, 'h10712, 'h10722, 'h10a60, 'h21f8e, 'h21f8f, 'h21f8d, 'h10732, 'h10742, 'h10a61, 'h10752, 'h10762, 'h10a62, 'h10772, 'h10782, 'h10a63, 'h10792, 'h10c62, 'h107a2, 'h10a64, 'h107b2, 'h103bc, 'h107c2, 'h10a65, 'h107d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e2, 'h10a66, 'h107f2, 'h10802, 'h10a67, 'h10812, 'h10822, 'h10a68, 'h10832, 'h10842, 'h10a69, 'h10c62, 'h10852, 'h10862, 'h10a6a, 'h103bc, 'h10872, 'h10882, 'h10a6b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10892, 'h108a2, 'h10a6c, 'h108b2, 'h108c2, 'h10a6d, 'h108d2, 'h106e2, 'h10a6e, 'h10c72, 'h106f2, 'h10702, 'h10a6f, 'h10712, 'h103bc, 'h10722, 'h10a70, 'h10732, 'h21f8e, 'h21f8f, 'h21f8d, 'h10742, 'h10a71, 'h10752, 'h10762, 'h10a72, 'h10772, 'h10782, 'h10a73, 'h10792, 'h10c72, 'h107a2, 'h10a74, 'h107b2, 'h107c2, 'h10a75, 'h103bc, 'h107d2, 'h107e2, 'h10a76, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f2, 'h10802, 'h10a77, 'h10812, 'h10822, 'h10a78, 'h10832, 'h10842, 'h10a79, 'h10c72, 'h10852, 'h10862, 'h10a7a, 'h10872, 'h103bc, 'h10882, 'h10a7b, 'h10892, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a2, 'h10a7c, 'h108b2, 'h108c2, 'h10a7d, 'h108d2, 'h106e2, 'h10a7e, 'h10c82, 'h106f2, 'h10702, 'h10a7f, 'h10712, 'h10722, 'h10a80, 'h103bc, 'h10732, 'h10742, 'h10a81, 'h21f8e, 'h21f8f, 'h21f8d, 'h10752, 'h10762, 'h10a82, 'h10772, 'h10782, 'h10a83, 'h10792, 'h10c82, 'h107a2, 'h10a84, 'h107b2, 'h107c2, 'h10a85, 'h107d2, 'h103bc, 'h107e2, 'h10a86, 'h107f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10802, 'h10a87, 'h10812, 'h10822, 'h10a88, 'h10832, 'h10842, 'h10a89, 'h10c82, 'h10852, 'h10862, 'h10a8a, 'h10872, 'h10882, 'h10a8b, 'h103bc, 'h10892, 'h108a2, 'h10a8c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b2, 'h108c2, 'h10a8d, 'h108d2, 'h106e2, 'h10a8e, 'h10c92, 'h106f2, 'h10702, 'h10a8f, 'h10712, 'h10722, 'h10a90, 'h10732, 'h103bc, 'h10742, 'h10a91, 'h10752, 'h21f8e, 'h21f8f, 'h21f8d, 'h10762, 'h10a92, 'h10772, 'h10782, 'h10a93, 'h10792, 'h10c92, 'h107a2, 'h10a94, 'h107b2, 'h107c2, 'h10a95, 'h107d2, 'h107e2, 'h10a96, 'h103bc, 'h107f2, 'h10802, 'h10a97, 'h21f8e, 'h21f8f, 'h21f8d, 'h10812, 'h10822, 'h10a98, 'h10832, 'h10842, 'h10a99, 'h10c92, 'h10852, 'h10862, 'h10a9a, 'h10872, 'h10882, 'h10a9b, 'h10892, 'h103bc, 'h108a2, 'h10a9c, 'h108b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c2, 'h10a9d, 'h108d2, 'h106e2, 'h10a9e, 'h10ca2, 'h106f2, 'h10702, 'h10a9f, 'h10712, 'h10722, 'h10aa0, 'h10732, 'h10742, 'h10aa1, 'h103bc, 'h10752, 'h10762, 'h10aa2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10772, 'h10782, 'h10aa3, 'h10792, 'h10ca2, 'h107a2, 'h10aa4, 'h107b2, 'h107c2, 'h10aa5, 'h107d2, 'h107e2, 'h10aa6, 'h107f2, 'h103bc, 'h10802, 'h10aa7, 'h10812, 'h21f8e, 'h21f8f, 'h21f8d, 'h10822, 'h10aa8, 'h10832, 'h10842, 'h10aa9, 'h10ca2, 'h10852, 'h10862, 'h10aaa, 'h10872, 'h10882, 'h10aab, 'h10892, 'h108a2, 'h10aac, 'h103bc, 'h108b2, 'h108c2, 'h10aad, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d2, 'h106e2, 'h10aae, 'h10cb2, 'h106f2, 'h10702, 'h10aaf, 'h10712, 'h10722, 'h10ab0, 'h10732, 'h10742, 'h10ab1, 'h10752, 'h103bc, 'h10762, 'h10ab2, 'h10772, 'h21f8e, 'h21f8f, 'h21f8d, 'h10782, 'h10ab3, 'h10792, 'h10cb2, 'h107a2, 'h10ab4, 'h107b2, 'h107c2, 'h10ab5, 'h107d2, 'h107e2, 'h10ab6, 'h107f2, 'h10802, 'h10ab7, 'h103bc, 'h10812, 'h10822, 'h10ab8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10832, 'h10842, 'h10ab9, 'h10cb2, 'h10852, 'h10862, 'h10aba, 'h10872, 'h10882, 'h10abb, 'h10892, 'h108a2, 'h10abc, 'h108b2, 'h103bc, 'h108c2, 'h10abd, 'h108d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h10abe, 'h10cc2, 'h106f2, 'h10702, 'h10abf, 'h10712, 'h10722, 'h10ac0, 'h10732, 'h10742, 'h10ac1, 'h10752, 'h10762, 'h10ac2, 'h103bc, 'h10772, 'h10782, 'h10ac3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10792, 'h10cc2, 'h107a2, 'h10ac4, 'h107b2, 'h107c2, 'h10ac5, 'h107d2, 'h107e2, 'h10ac6, 'h107f2, 'h10802, 'h10ac7, 'h10812, 'h103bc, 'h10822, 'h10ac8, 'h10832, 'h21f8e, 'h21f8f, 'h21f8d, 'h10842, 'h10ac9, 'h10cc2, 'h10852, 'h10862, 'h10aca, 'h10872, 'h10882, 'h10acb, 'h10892, 'h108a2, 'h10acc, 'h108b2, 'h108c2, 'h10acd, 'h103bc, 'h108d2, 'h106e2, 'h10ace, 'h10cd2, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f2, 'h10702, 'h10acf, 'h10712, 'h10722, 'h10ad0, 'h10732, 'h10742, 'h10ad1, 'h10752, 'h10762, 'h10ad2, 'h10772, 'h103bc, 'h10782, 'h10ad3, 'h10792, 'h10cd2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a2, 'h10ad4, 'h107b2, 'h107c2, 'h10ad5, 'h107d2, 'h107e2, 'h10ad6, 'h107f2, 'h10802, 'h10ad7, 'h10812, 'h10822, 'h10ad8, 'h103bc, 'h10832, 'h10842, 'h10ad9, 'h10cd2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10852, 'h10862, 'h10ada, 'h10872, 'h10882, 'h10adb, 'h10892, 'h108a2, 'h10adc, 'h108b2, 'h108c2, 'h10add, 'h108d2, 'h103bc, 'h106e2, 'h108de, 'h10ae2, 'h106f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10702, 'h108df, 'h10712, 'h10722, 'h108e0, 'h10732, 'h10742, 'h108e1, 'h10752, 'h10762, 'h108e2, 'h10772, 'h10782, 'h108e3, 'h103bc, 'h10792, 'h10ae2, 'h107a2, 'h108e4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b2, 'h107c2, 'h108e5, 'h107d2, 'h107e2, 'h108e6, 'h107f2, 'h10802, 'h108e7, 'h10812, 'h10822, 'h108e8, 'h10832, 'h103bc, 'h10842, 'h108e9, 'h10ae2, 'h10852, 'h21f8e, 'h21f8f, 'h21f8d, 'h10862, 'h108ea, 'h10872, 'h10882, 'h108eb, 'h10892, 'h108a2, 'h108ec, 'h108b2, 'h108c2, 'h108ed, 'h108d2, 'h106e2, 'h108ee, 'h10af2, 'h103bc, 'h106f2, 'h10702, 'h108ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h10712, 'h10722, 'h108f0, 'h10732, 'h10742, 'h108f1, 'h10752, 'h10762, 'h108f2, 'h10772, 'h10782, 'h108f3, 'h10792, 'h10af2, 'h103bc, 'h107a2, 'h108f4, 'h107b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c2, 'h108f5, 'h107d2, 'h107e2, 'h108f6, 'h107f2, 'h10802, 'h108f7, 'h10812, 'h10822, 'h108f8, 'h10832, 'h10842, 'h108f9, 'h10af2, 'h103bc, 'h10852, 'h10862, 'h108fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h10872, 'h10882, 'h108fb, 'h10892, 'h108a2, 'h108fc, 'h108b2, 'h108c2, 'h108fd, 'h108d2, 'h106e2, 'h108fe, 'h10b02, 'h106f2, 'h103bc, 'h10702, 'h108ff, 'h10712, 'h21f8e, 'h21f8f, 'h21f8d, 'h10722, 'h10900, 'h10732, 'h10742, 'h10901, 'h10752, 'h10762, 'h10902, 'h10772, 'h10782, 'h10903, 'h10792, 'h10b02, 'h107a2, 'h10904, 'h103bc, 'h107b2, 'h107c2, 'h10905, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d2, 'h107e2, 'h10906, 'h107f2, 'h10802, 'h10907, 'h10812, 'h10822, 'h10908, 'h10832, 'h10842, 'h10909, 'h10b02, 'h10852, 'h103bc, 'h10862, 'h1090a, 'h10872, 'h21f8e, 'h21f8f, 'h21f8d, 'h10882, 'h1090b, 'h10892, 'h108a2, 'h1090c, 'h108b2, 'h108c2, 'h1090d, 'h108d2, 'h106e2, 'h1090e, 'h10b12, 'h106f2, 'h10702, 'h1090f, 'h103bc, 'h10712, 'h10722, 'h10910, 'h21f8e, 'h21f8f, 'h21f8d, 'h10732, 'h10742, 'h10911, 'h10752, 'h10762, 'h10912, 'h10772, 'h10782, 'h10913, 'h10792, 'h10b12, 'h107a2, 'h10914, 'h107b2, 'h103bc, 'h107c2, 'h10915, 'h107d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e2, 'h10916, 'h107f2, 'h10802, 'h10917, 'h10812, 'h10822, 'h10918, 'h10832, 'h10842, 'h10919, 'h10b12, 'h10852, 'h10862, 'h1091a, 'h103bc, 'h10872, 'h10882, 'h1091b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10892, 'h108a2, 'h1091c, 'h108b2, 'h108c2, 'h1091d, 'h108d2, 'h106e2, 'h1091e, 'h10b22, 'h106f2, 'h10702, 'h1091f, 'h10712, 'h103bc, 'h10722, 'h10920, 'h10732, 'h21f8e, 'h21f8f, 'h21f8d, 'h10742, 'h10921, 'h10752, 'h10762, 'h10922, 'h10772, 'h10782, 'h10923, 'h10792, 'h10b22, 'h107a2, 'h10924, 'h107b2, 'h107c2, 'h10925, 'h103bc, 'h107d2, 'h107e2, 'h10926, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f2, 'h10802, 'h10927, 'h10812, 'h10822, 'h10928, 'h10832, 'h10842, 'h10929, 'h10b22, 'h10852, 'h10862, 'h1092a, 'h10872, 'h103bc, 'h10882, 'h1092b, 'h10892, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a2, 'h1092c, 'h108b2, 'h108c2, 'h1092d, 'h108d2, 'h106e2, 'h1092e, 'h10b32, 'h106f2, 'h10702, 'h1092f, 'h10712, 'h10722, 'h10930, 'h103bc, 'h10732, 'h10742, 'h10931, 'h21f8e, 'h21f8f, 'h21f8d, 'h10752, 'h10762, 'h10932, 'h10772, 'h10782, 'h10933, 'h10792, 'h10b32, 'h107a2, 'h10934, 'h107b2, 'h107c2, 'h10935, 'h107d2, 'h103bc, 'h107e2, 'h10936, 'h107f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10802, 'h10937, 'h10812, 'h10822, 'h10938, 'h10832, 'h10842, 'h10939, 'h10b32, 'h10852, 'h10862, 'h1093a, 'h10872, 'h10882, 'h1093b, 'h103bc, 'h10892, 'h108a2, 'h1093c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b2, 'h108c2, 'h1093d, 'h108d2, 'h106e2, 'h1093e, 'h10b42, 'h106f2, 'h10702, 'h1093f, 'h10712, 'h10722, 'h10940, 'h10732, 'h103bc, 'h10742, 'h10941, 'h10752, 'h21f8e, 'h21f8f, 'h21f8d, 'h10762, 'h10942, 'h10772, 'h10782, 'h10943, 'h10792, 'h10b42, 'h107a2, 'h10944, 'h107b2, 'h107c2, 'h10945, 'h107d2, 'h107e2, 'h10946, 'h103bc, 'h107f2, 'h10802, 'h10947, 'h21f8e, 'h21f8f, 'h21f8d, 'h10812, 'h10822, 'h10948, 'h10832, 'h10842, 'h10949, 'h10b42, 'h10852, 'h10862, 'h1094a, 'h10872, 'h10882, 'h1094b, 'h10892, 'h103bc, 'h108a2, 'h1094c, 'h108b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c2, 'h1094d, 'h108d2, 'h106e2, 'h1094e, 'h10b52, 'h106f2, 'h10702, 'h1094f, 'h10712, 'h10722, 'h10950, 'h10732, 'h10742, 'h10951, 'h103bc, 'h10752, 'h10762, 'h10952, 'h21f8e, 'h21f8f, 'h21f8d, 'h10772, 'h10782, 'h10953, 'h10792, 'h10b52, 'h107a2, 'h10954, 'h107b2, 'h107c2, 'h10955, 'h107d2, 'h107e2, 'h10956, 'h107f2, 'h103bc, 'h10802, 'h10957, 'h10812, 'h21f8e, 'h21f8f, 'h21f8d, 'h10822, 'h10958, 'h10832, 'h10842, 'h10959, 'h10b52, 'h10852, 'h10862, 'h1095a, 'h10872, 'h10882, 'h1095b, 'h10892, 'h108a2, 'h1095c, 'h103bc, 'h108b2, 'h108c2, 'h1095d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d2, 'h106e2, 'h1095e, 'h10b62, 'h106f2, 'h10702, 'h1095f, 'h10712, 'h10722, 'h10960, 'h10732, 'h10742, 'h10961, 'h10752, 'h103bc, 'h10762, 'h10962, 'h10772, 'h21f8e, 'h21f8f, 'h21f8d, 'h10782, 'h10963, 'h10792, 'h10b62, 'h107a2, 'h10964, 'h107b2, 'h107c2, 'h10965, 'h107d2, 'h107e2, 'h10966, 'h107f2, 'h10802, 'h10967, 'h103bc, 'h10812, 'h10822, 'h10968, 'h21f8e, 'h21f8f, 'h21f8d, 'h10832, 'h10842, 'h10969, 'h10b62, 'h10852, 'h10862, 'h1096a, 'h10872, 'h10882, 'h1096b, 'h10892, 'h108a2, 'h1096c, 'h108b2, 'h103bc, 'h108c2, 'h1096d, 'h108d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1096e, 'h10b72, 'h106f2, 'h10702, 'h1096f, 'h10712, 'h10722, 'h10970, 'h10732, 'h10742, 'h10971, 'h10752, 'h10762, 'h10972, 'h103bc, 'h10772, 'h10782, 'h10973, 'h21f8e, 'h21f8f, 'h21f8d, 'h10792, 'h10b72, 'h107a2, 'h10974, 'h107b2, 'h107c2, 'h10975, 'h107d2, 'h107e2, 'h10976, 'h107f2, 'h10802, 'h10977, 'h10812, 'h103bc, 'h10822, 'h10978, 'h10832, 'h21f8e, 'h21f8f, 'h21f8d, 'h10842, 'h10979, 'h10b72, 'h10852, 'h10862, 'h1097a, 'h10872, 'h10882, 'h1097b, 'h10892, 'h108a2, 'h1097c, 'h108b2, 'h108c2, 'h1097d, 'h103bc, 'h108d2, 'h106e2, 'h1097e, 'h10b82, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f2, 'h10702, 'h1097f, 'h10712, 'h10722, 'h10980, 'h10732, 'h10742, 'h10981, 'h10752, 'h10762, 'h10982, 'h10772, 'h103bc, 'h10782, 'h10983, 'h10792, 'h10b82, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a2, 'h10984, 'h107b2, 'h107c2, 'h10985, 'h107d2, 'h107e2, 'h10986, 'h107f2, 'h10802, 'h10987, 'h10812, 'h10822, 'h10988, 'h103bc, 'h10832, 'h10842, 'h10989, 'h10b82, 'h21f8e, 'h21f8f, 'h21f8d, 'h10852, 'h10862, 'h1098a, 'h10872, 'h10882, 'h1098b, 'h10892, 'h108a2, 'h1098c, 'h108b2, 'h108c2, 'h1098d, 'h108d2, 'h103bc, 'h106e2, 'h1098e, 'h10b92, 'h106f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10702, 'h1098f, 'h10712, 'h10722, 'h10990, 'h10732, 'h10742, 'h10991, 'h10752, 'h10762, 'h10992, 'h10772, 'h10782, 'h10993, 'h103bc, 'h10792, 'h10b92, 'h107a2, 'h10994, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b2, 'h107c2, 'h10995, 'h107d2, 'h107e2, 'h10996, 'h107f2, 'h10802, 'h10997, 'h10812, 'h10822, 'h10998, 'h10832, 'h103bc, 'h10842, 'h10999, 'h10b92, 'h10852, 'h21f8e, 'h21f8f, 'h21f8d, 'h10862, 'h1099a, 'h10872, 'h10882, 'h1099b, 'h10892, 'h108a2, 'h1099c, 'h108b2, 'h108c2, 'h1099d, 'h108d2, 'h106e2, 'h1099e, 'h10ba2, 'h103bc, 'h106f2, 'h10702, 'h1099f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10712, 'h10722, 'h109a0, 'h10732, 'h10742, 'h109a1, 'h10752, 'h10762, 'h109a2, 'h10772, 'h10782, 'h109a3, 'h10792, 'h10ba2, 'h103bc, 'h107a2, 'h109a4, 'h107b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c2, 'h109a5, 'h107d2, 'h107e2, 'h109a6, 'h107f2, 'h10802, 'h109a7, 'h10812, 'h10822, 'h109a8, 'h10832, 'h10842, 'h109a9, 'h10ba2, 'h103bc, 'h10852, 'h10862, 'h109aa, 'h21f8e, 'h21f8f, 'h21f8d, 'h10872, 'h10882, 'h109ab, 'h10892, 'h108a2, 'h109ac, 'h108b2, 'h108c2, 'h109ad, 'h108d2, 'h106e2, 'h109ae, 'h10bb2, 'h106f2, 'h103bc, 'h10702, 'h109af, 'h10712, 'h21f8e, 'h21f8f, 'h21f8d, 'h10722, 'h109b0, 'h10732, 'h10742, 'h109b1, 'h10752, 'h10762, 'h109b2, 'h10772, 'h10782, 'h109b3, 'h10792, 'h10bb2, 'h107a2, 'h109b4, 'h103bc, 'h107b2, 'h107c2, 'h109b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d2, 'h107e2, 'h109b6, 'h107f2, 'h10802, 'h109b7, 'h10812, 'h10822, 'h109b8, 'h10832, 'h10842, 'h109b9, 'h10bb2, 'h10852, 'h103bc, 'h10862, 'h109ba, 'h10872, 'h21f8e, 'h21f8f, 'h21f8d, 'h10882, 'h109bb, 'h10892, 'h108a2, 'h109bc, 'h108b2, 'h108c2, 'h109bd, 'h108d2, 'h106e2, 'h109be, 'h10bc2, 'h106f2, 'h10702, 'h109bf, 'h103bc, 'h10712, 'h10722, 'h109c0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10732, 'h10742, 'h109c1, 'h10752, 'h10762, 'h109c2, 'h10772, 'h10782, 'h109c3, 'h10792, 'h10bc2, 'h107a2, 'h109c4, 'h107b2, 'h103bc, 'h107c2, 'h109c5, 'h107d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e2, 'h109c6, 'h107f2, 'h10802, 'h109c7, 'h10812, 'h10822, 'h109c8, 'h10832, 'h10842, 'h109c9, 'h10bc2, 'h10852, 'h10862, 'h109ca, 'h103bc, 'h10872, 'h10882, 'h109cb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10892, 'h108a2, 'h109cc, 'h108b2, 'h108c2, 'h109cd, 'h108d2, 'h106e2, 'h109ce, 'h10bd2, 'h106f2, 'h10702, 'h109cf, 'h10712, 'h103bc, 'h10722, 'h109d0, 'h10732, 'h21f8e, 'h21f8f, 'h21f8d, 'h10742, 'h109d1, 'h10752, 'h10762, 'h109d2, 'h10772, 'h10782, 'h109d3, 'h10792, 'h10bd2, 'h107a2, 'h109d4, 'h107b2, 'h107c2, 'h109d5, 'h103bc, 'h107d2, 'h107e2, 'h109d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f2, 'h10802, 'h109d7, 'h10812, 'h10822, 'h109d8, 'h10832, 'h10842, 'h109d9, 'h10bd2, 'h10852, 'h10862, 'h109da, 'h10872, 'h103bc, 'h10882, 'h109db, 'h10892, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a2, 'h109dc, 'h108b2, 'h108c2, 'h109dd, 'h108d2, 'h106e2, 'h109de, 'h10be2, 'h106f2, 'h10702, 'h109df, 'h10712, 'h10722, 'h109e0, 'h103bc, 'h10732, 'h10742, 'h109e1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10752, 'h10762, 'h109e2, 'h10772, 'h10782, 'h109e3, 'h10792, 'h10be2, 'h107a2, 'h109e4, 'h107b2, 'h107c2, 'h109e5, 'h107d2, 'h103bc, 'h107e2, 'h109e6, 'h107f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10802, 'h109e7, 'h10812, 'h10822, 'h109e8, 'h10832, 'h10842, 'h109e9, 'h10be2, 'h10852, 'h10862, 'h109ea, 'h10872, 'h10882, 'h109eb, 'h103bc, 'h10892, 'h108a2, 'h109ec, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b2, 'h108c2, 'h109ed, 'h108d2, 'h106e2, 'h109ee, 'h10bf2, 'h106f2, 'h10702, 'h109ef, 'h10712, 'h10722, 'h109f0, 'h10732, 'h103bc, 'h10742, 'h109f1, 'h10752, 'h21f8e, 'h21f8f, 'h21f8d, 'h10762, 'h109f2, 'h10772, 'h10782, 'h109f3, 'h10792, 'h10bf2, 'h107a2, 'h109f4, 'h107b2, 'h107c2, 'h109f5, 'h107d2, 'h107e2, 'h109f6, 'h103bc, 'h107f2, 'h10802, 'h109f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10812, 'h10822, 'h109f8, 'h10832, 'h10842, 'h109f9, 'h10bf2, 'h10852, 'h10862, 'h109fa, 'h10872, 'h10882, 'h109fb, 'h10892, 'h103bc, 'h108a2, 'h109fc, 'h108b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c2, 'h109fd, 'h108d2, 'h106e2, 'h109fe, 'h10c02, 'h106f2, 'h10702, 'h109ff, 'h10712, 'h10722, 'h10a00, 'h10732, 'h10742, 'h10a01, 'h103bc, 'h10752, 'h10762, 'h10a02, 'h21f8e, 'h21f8f, 'h21f8d, 'h10772, 'h10782, 'h10a03, 'h10792, 'h10c02, 'h107a2, 'h10a04, 'h107b2, 'h107c2, 'h10a05, 'h107d2, 'h107e2, 'h10a06, 'h107f2, 'h103bc, 'h10802, 'h10a07, 'h10812, 'h21f8e, 'h21f8f, 'h21f8d, 'h10822, 'h10a08, 'h10832, 'h10842, 'h10a09, 'h10c02, 'h10852, 'h10862, 'h10a0a, 'h10872, 'h10882, 'h10a0b, 'h10892, 'h108a2, 'h10a0c, 'h103bc, 'h108b2, 'h108c2, 'h10a0d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d2, 'h106e2, 'h10a0e, 'h10c12, 'h106f2, 'h10702, 'h10a0f, 'h10712, 'h10722, 'h10a10, 'h10732, 'h10742, 'h10a11, 'h10752, 'h103bc, 'h10762, 'h10a12, 'h10772, 'h21f8e, 'h21f8f, 'h21f8d, 'h10782, 'h10a13, 'h10792, 'h10c12, 'h107a2, 'h10a14, 'h107b2, 'h107c2, 'h10a15, 'h107d2, 'h107e2, 'h10a16, 'h107f2, 'h10802, 'h10a17, 'h103bc, 'h10812, 'h10822, 'h10a18, 'h21f8e, 'h21f8f, 'h21f8d, 'h10832, 'h10842, 'h10a19, 'h10c12, 'h10852, 'h10862, 'h10a1a, 'h10872, 'h10882, 'h10a1b, 'h10892, 'h108a2, 'h10a1c, 'h108b2, 'h103bc, 'h108c2, 'h10a1d, 'h108d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h10a1e, 'h10c22, 'h106f2, 'h10702, 'h10a1f, 'h10712, 'h10722, 'h10a20, 'h10732, 'h10742, 'h10a21, 'h10752, 'h10762, 'h10a22, 'h103bc, 'h10772, 'h10782, 'h10a23, 'h21f8e, 'h21f8f, 'h21f8d, 'h10792, 'h10c22, 'h107a2, 'h10a24, 'h107b2, 'h107c2, 'h10a25, 'h107d2, 'h107e2, 'h10a26, 'h107f2, 'h10802, 'h10a27, 'h10812, 'h103bc, 'h10822, 'h10a28, 'h10832, 'h21f8e, 'h21f8f, 'h21f8d, 'h10842, 'h10a29, 'h10c22, 'h10852, 'h10862, 'h10a2a, 'h10872, 'h10882, 'h10a2b, 'h10892, 'h108a2, 'h10a2c, 'h108b2, 'h108c2, 'h10a2d, 'h103bc, 'h108d2, 'h106e2, 'h10a2e, 'h10c32, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f2, 'h10702, 'h10a2f, 'h10712, 'h10722, 'h10a30, 'h10732, 'h10742, 'h10a31, 'h10752, 'h10762, 'h10a32, 'h10772, 'h103bc, 'h10782, 'h10a33, 'h10792, 'h10c32, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a2, 'h10a34, 'h107b2, 'h107c2, 'h10a35, 'h107d2, 'h107e2, 'h10a36, 'h107f2, 'h10802, 'h10a37, 'h10812, 'h10822, 'h10a38, 'h103bc, 'h10832, 'h10842, 'h10a39, 'h10c32, 'h21f8e, 'h21f8f, 'h21f8d, 'h10852, 'h10862, 'h10a3a, 'h10872, 'h10882, 'h10a3b, 'h10892, 'h108a2, 'h10a3c, 'h108b2, 'h108c2, 'h10a3d, 'h108d2, 'h103bc, 'h106e2, 'h10a3e, 'h10c42, 'h106f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10702, 'h10a3f, 'h10712, 'h10722, 'h10a40, 'h10732, 'h10742, 'h10a41, 'h10752, 'h10762, 'h10a42, 'h10772, 'h10782, 'h10a43, 'h103bc, 'h10792, 'h10c42, 'h107a2, 'h10a44, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b2, 'h107c2, 'h10a45, 'h107d2, 'h107e2, 'h10a46, 'h107f2, 'h10802, 'h10a47, 'h10812, 'h10822, 'h10a48, 'h10832, 'h103bc, 'h10842, 'h10a49, 'h10c42, 'h10852, 'h21f8e, 'h21f8f, 'h21f8d, 'h10862, 'h10a4a, 'h10872, 'h10882, 'h10a4b, 'h10892, 'h108a2, 'h10a4c, 'h108b2, 'h108c2, 'h10a4d, 'h108d2, 'h106e2, 'h10a4e, 'h10c52, 'h103bc, 'h106f2, 'h10702, 'h10a4f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10712, 'h10722, 'h10a50, 'h10732, 'h10742, 'h10a51, 'h10752, 'h10762, 'h10a52, 'h10772, 'h10782, 'h10a53, 'h10792, 'h10c52, 'h103bc, 'h107a2, 'h10a54, 'h107b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c2, 'h10a55, 'h107d2, 'h107e2, 'h10a56, 'h107f2, 'h10802, 'h10a57, 'h10812, 'h10822, 'h10a58, 'h10832, 'h10842, 'h10a59, 'h10c52, 'h103bc, 'h10852, 'h10862, 'h10a5a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10872, 'h10882, 'h10a5b, 'h10892, 'h108a2, 'h10a5c, 'h108b2, 'h108c2, 'h10a5d, 'h108d2, 'h106e2, 'h10a5e, 'h10c62, 'h106f2, 'h103bc, 'h10702, 'h10a5f, 'h10712, 'h21f8e, 'h21f8f, 'h21f8d, 'h10722, 'h10a60, 'h10732, 'h10742, 'h10a61, 'h10752, 'h10762, 'h10a62, 'h10772, 'h10782, 'h10a63, 'h10792, 'h10c62, 'h107a2, 'h10a64, 'h103bc, 'h107b2, 'h107c2, 'h10a65, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d2, 'h107e2, 'h10a66, 'h107f2, 'h10802, 'h10a67, 'h10812, 'h10822, 'h10a68, 'h10832, 'h10842, 'h10a69, 'h10c62, 'h10852, 'h103bc, 'h10862, 'h10a6a, 'h10872, 'h21f8e, 'h21f8f, 'h21f8d, 'h10882, 'h10a6b, 'h10892, 'h108a2, 'h10a6c, 'h108b2, 'h108c2, 'h10a6d, 'h108d2, 'h106e2, 'h10a6e, 'h10c72, 'h106f2, 'h10702, 'h10a6f, 'h103bc, 'h10712, 'h10722, 'h10a70, 'h21f8e, 'h21f8f, 'h21f8d, 'h10732, 'h10742, 'h10a71, 'h10752, 'h10762, 'h10a72, 'h10772, 'h10782, 'h10a73, 'h10792, 'h10c72, 'h107a2, 'h10a74, 'h107b2, 'h103bc, 'h107c2, 'h10a75, 'h107d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e2, 'h10a76, 'h107f2, 'h10802, 'h10a77, 'h10812, 'h10822, 'h10a78, 'h10832, 'h10842, 'h10a79, 'h10c72, 'h10852, 'h10862, 'h10a7a, 'h103bc, 'h10872, 'h10882, 'h10a7b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10892, 'h108a2, 'h10a7c, 'h108b2, 'h108c2, 'h10a7d, 'h108d2, 'h106e2, 'h10a7e, 'h10c82, 'h106f2, 'h10702, 'h10a7f, 'h10712, 'h103bc, 'h10722, 'h10a80, 'h10732, 'h21f8e, 'h21f8f, 'h21f8d, 'h10742, 'h10a81, 'h10752, 'h10762, 'h10a82, 'h10772, 'h10782, 'h10a83, 'h10792, 'h10c82, 'h107a2, 'h10a84, 'h107b2, 'h107c2, 'h10a85, 'h103bc, 'h107d2, 'h107e2, 'h10a86, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f2, 'h10802, 'h10a87, 'h10812, 'h10822, 'h10a88, 'h10832, 'h10842, 'h10a89, 'h10c82, 'h10852, 'h10862, 'h10a8a, 'h10872, 'h103bc, 'h10882, 'h10a8b, 'h10892, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a2, 'h10a8c, 'h108b2, 'h108c2, 'h10a8d, 'h108d2, 'h106e2, 'h10a8e, 'h10c92, 'h106f2, 'h10702, 'h10a8f, 'h10712, 'h10722, 'h10a90, 'h103bc, 'h10732, 'h10742, 'h10a91, 'h21f8e, 'h21f8f, 'h21f8d, 'h10752, 'h10762, 'h10a92, 'h10772, 'h10782, 'h10a93, 'h10792, 'h10c92, 'h107a2, 'h10a94, 'h107b2, 'h107c2, 'h10a95, 'h107d2, 'h103bc, 'h107e2, 'h10a96, 'h107f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10802, 'h10a97, 'h10812, 'h10822, 'h10a98, 'h10832, 'h10842, 'h10a99, 'h10c92, 'h10852, 'h10862, 'h10a9a, 'h10872, 'h10882, 'h10a9b, 'h103bc, 'h10892, 'h108a2, 'h10a9c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b2, 'h108c2, 'h10a9d, 'h108d2, 'h106e2, 'h10a9e, 'h10ca2, 'h106f2, 'h10702, 'h10a9f, 'h10712, 'h10722, 'h10aa0, 'h10732, 'h103bc, 'h10742, 'h10aa1, 'h10752, 'h21f8e, 'h21f8f, 'h21f8d, 'h10762, 'h10aa2, 'h10772, 'h10782, 'h10aa3, 'h10792, 'h10ca2, 'h107a2, 'h10aa4, 'h107b2, 'h107c2, 'h10aa5, 'h107d2, 'h107e2, 'h10aa6, 'h103bc, 'h107f2, 'h10802, 'h10aa7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10812, 'h10822, 'h10aa8, 'h10832, 'h10842, 'h10aa9, 'h10ca2, 'h10852, 'h10862, 'h10aaa, 'h10872, 'h10882, 'h10aab, 'h10892, 'h103bc, 'h108a2, 'h10aac, 'h108b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c2, 'h10aad, 'h108d2, 'h106e2, 'h10aae, 'h10cb2, 'h106f2, 'h10702, 'h10aaf, 'h10712, 'h10722, 'h10ab0, 'h10732, 'h10742, 'h10ab1, 'h103bc, 'h10752, 'h10762, 'h10ab2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10772, 'h10782, 'h10ab3, 'h10792, 'h10cb2, 'h107a2, 'h10ab4, 'h107b2, 'h107c2, 'h10ab5, 'h107d2, 'h107e2, 'h10ab6, 'h107f2, 'h103bc, 'h10802, 'h10ab7, 'h10812, 'h21f8e, 'h21f8f, 'h21f8d, 'h10822, 'h10ab8, 'h10832, 'h10842, 'h10ab9, 'h10cb2, 'h10852, 'h10862, 'h10aba, 'h10872, 'h10882, 'h10abb, 'h10892, 'h108a2, 'h10abc, 'h103bc, 'h108b2, 'h108c2, 'h10abd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d2, 'h106e2, 'h10abe, 'h10cc2, 'h106f2, 'h10702, 'h10abf, 'h10712, 'h10722, 'h10ac0, 'h10732, 'h10742, 'h10ac1, 'h10752, 'h103bc, 'h10762, 'h10ac2, 'h10772, 'h21f8e, 'h21f8f, 'h21f8d, 'h10782, 'h10ac3, 'h10792, 'h10cc2, 'h107a2, 'h10ac4, 'h107b2, 'h107c2, 'h10ac5, 'h107d2, 'h107e2, 'h10ac6, 'h107f2, 'h10802, 'h10ac7, 'h103bc, 'h10812, 'h10822, 'h10ac8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10832, 'h10842, 'h10ac9, 'h10cc2, 'h10852, 'h10862, 'h10aca, 'h10872, 'h10882, 'h10acb, 'h10892, 'h108a2, 'h10acc, 'h108b2, 'h103bc, 'h108c2, 'h10acd, 'h108d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h10ace, 'h10cd2, 'h106f2, 'h10702, 'h10acf, 'h10712, 'h10722, 'h10ad0, 'h10732, 'h10742, 'h10ad1, 'h10752, 'h10762, 'h10ad2, 'h103bc, 'h10772, 'h10782, 'h10ad3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10792, 'h10cd2, 'h107a2, 'h10ad4, 'h107b2, 'h107c2, 'h10ad5, 'h107d2, 'h107e2, 'h10ad6, 'h107f2, 'h10802, 'h10ad7, 'h10812, 'h103bc, 'h10822, 'h10ad8, 'h10832, 'h21f8e, 'h21f8f, 'h21f8d, 'h10842, 'h10ad9, 'h10cd2, 'h10852, 'h10862, 'h10ada, 'h10872, 'h10882, 'h10adb, 'h10892, 'h108a2, 'h10adc, 'h108b2, 'h108c2, 'h10add, 'h103bc, 'h108d2, 'h106e3, 'h108de, 'h10ae3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f3, 'h10703, 'h108df, 'h10713, 'h10723, 'h108e0, 'h10733, 'h10743, 'h108e1, 'h10753, 'h10763, 'h108e2, 'h10773, 'h103bc, 'h10783, 'h108e3, 'h10793, 'h10ae3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a3, 'h108e4, 'h107b3, 'h107c3, 'h108e5, 'h107d3, 'h107e3, 'h108e6, 'h107f3, 'h10803, 'h108e7, 'h10813, 'h10823, 'h108e8, 'h103bc, 'h10833, 'h10843, 'h108e9, 'h10ae3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10853, 'h10863, 'h108ea, 'h10873, 'h10883, 'h108eb, 'h10893, 'h108a3, 'h108ec, 'h108b3, 'h108c3, 'h108ed, 'h108d3, 'h103bc, 'h106e3, 'h108ee, 'h10af3, 'h106f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10703, 'h108ef, 'h10713, 'h10723, 'h108f0, 'h10733, 'h10743, 'h108f1, 'h10753, 'h10763, 'h108f2, 'h10773, 'h10783, 'h108f3, 'h103bc, 'h10793, 'h10af3, 'h107a3, 'h108f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b3, 'h107c3, 'h108f5, 'h107d3, 'h107e3, 'h108f6, 'h107f3, 'h10803, 'h108f7, 'h10813, 'h10823, 'h108f8, 'h10833, 'h103bc, 'h10843, 'h108f9, 'h10af3, 'h10853, 'h21f8e, 'h21f8f, 'h21f8d, 'h10863, 'h108fa, 'h10873, 'h10883, 'h108fb, 'h10893, 'h108a3, 'h108fc, 'h108b3, 'h108c3, 'h108fd, 'h108d3, 'h106e3, 'h108fe, 'h10b03, 'h103bc, 'h106f3, 'h10703, 'h108ff, 'h21f8e, 'h21f8f, 'h21f8d, 'h10713, 'h10723, 'h10900, 'h10733, 'h10743, 'h10901, 'h10753, 'h10763, 'h10902, 'h10773, 'h10783, 'h10903, 'h10793, 'h10b03, 'h103bc, 'h107a3, 'h10904, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c3, 'h10905, 'h107d3, 'h107e3, 'h10906, 'h107f3, 'h10803, 'h10907, 'h10813, 'h10823, 'h10908, 'h10833, 'h10843, 'h10909, 'h10b03, 'h103bc, 'h10853, 'h10863, 'h1090a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10873, 'h10883, 'h1090b, 'h10893, 'h108a3, 'h1090c, 'h108b3, 'h108c3, 'h1090d, 'h108d3, 'h106e3, 'h1090e, 'h10b13, 'h106f3, 'h103bc, 'h10703, 'h1090f, 'h10713, 'h21f8e, 'h21f8f, 'h21f8d, 'h10723, 'h10910, 'h10733, 'h10743, 'h10911, 'h10753, 'h10763, 'h10912, 'h10773, 'h10783, 'h10913, 'h10793, 'h10b13, 'h107a3, 'h10914, 'h103bc, 'h107b3, 'h107c3, 'h10915, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d3, 'h107e3, 'h10916, 'h107f3, 'h10803, 'h10917, 'h10813, 'h10823, 'h10918, 'h10833, 'h10843, 'h10919, 'h10b13, 'h10853, 'h103bc, 'h10863, 'h1091a, 'h10873, 'h21f8e, 'h21f8f, 'h21f8d, 'h10883, 'h1091b, 'h10893, 'h108a3, 'h1091c, 'h108b3, 'h108c3, 'h1091d, 'h108d3, 'h106e3, 'h1091e, 'h10b23, 'h106f3, 'h10703, 'h1091f, 'h103bc, 'h10713, 'h10723, 'h10920, 'h21f8e, 'h21f8f, 'h21f8d, 'h10733, 'h10743, 'h10921, 'h10753, 'h10763, 'h10922, 'h10773, 'h10783, 'h10923, 'h10793, 'h10b23, 'h107a3, 'h10924, 'h107b3, 'h103bc, 'h107c3, 'h10925, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e3, 'h10926, 'h107f3, 'h10803, 'h10927, 'h10813, 'h10823, 'h10928, 'h10833, 'h10843, 'h10929, 'h10b23, 'h10853, 'h10863, 'h1092a, 'h103bc, 'h10873, 'h10883, 'h1092b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10893, 'h108a3, 'h1092c, 'h108b3, 'h108c3, 'h1092d, 'h108d3, 'h106e3, 'h1092e, 'h10b33, 'h106f3, 'h10703, 'h1092f, 'h10713, 'h103bc, 'h10723, 'h10930, 'h10733, 'h21f8e, 'h21f8f, 'h21f8d, 'h10743, 'h10931, 'h10753, 'h10763, 'h10932, 'h10773, 'h10783, 'h10933, 'h10793, 'h10b33, 'h107a3, 'h10934, 'h107b3, 'h107c3, 'h10935, 'h103bc, 'h107d3, 'h107e3, 'h10936, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f3, 'h10803, 'h10937, 'h10813, 'h10823, 'h10938, 'h10833, 'h10843, 'h10939, 'h10b33, 'h10853, 'h10863, 'h1093a, 'h10873, 'h103bc, 'h10883, 'h1093b, 'h10893, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a3, 'h1093c, 'h108b3, 'h108c3, 'h1093d, 'h108d3, 'h106e3, 'h1093e, 'h10b43, 'h106f3, 'h10703, 'h1093f, 'h10713, 'h10723, 'h10940, 'h103bc, 'h10733, 'h10743, 'h10941, 'h21f8e, 'h21f8f, 'h21f8d, 'h10753, 'h10763, 'h10942, 'h10773, 'h10783, 'h10943, 'h10793, 'h10b43, 'h107a3, 'h10944, 'h107b3, 'h107c3, 'h10945, 'h107d3, 'h103bc, 'h107e3, 'h10946, 'h107f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10803, 'h10947, 'h10813, 'h10823, 'h10948, 'h10833, 'h10843, 'h10949, 'h10b43, 'h10853, 'h10863, 'h1094a, 'h10873, 'h10883, 'h1094b, 'h103bc, 'h10893, 'h108a3, 'h1094c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b3, 'h108c3, 'h1094d, 'h108d3, 'h106e3, 'h1094e, 'h10b53, 'h106f3, 'h10703, 'h1094f, 'h10713, 'h10723, 'h10950, 'h10733, 'h103bc, 'h10743, 'h10951, 'h10753, 'h21f8e, 'h21f8f, 'h21f8d, 'h10763, 'h10952, 'h10773, 'h10783, 'h10953, 'h10793, 'h10b53, 'h107a3, 'h10954, 'h107b3, 'h107c3, 'h10955, 'h107d3, 'h107e3, 'h10956, 'h103bc, 'h107f3, 'h10803, 'h10957, 'h21f8e, 'h21f8f, 'h21f8d, 'h10813, 'h10823, 'h10958, 'h10833, 'h10843, 'h10959, 'h10b53, 'h10853, 'h10863, 'h1095a, 'h10873, 'h10883, 'h1095b, 'h10893, 'h103bc, 'h108a3, 'h1095c, 'h108b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c3, 'h1095d, 'h108d3, 'h106e3, 'h1095e, 'h10b63, 'h106f3, 'h10703, 'h1095f, 'h10713, 'h10723, 'h10960, 'h10733, 'h10743, 'h10961, 'h103bc, 'h10753, 'h10763, 'h10962, 'h21f8e, 'h21f8f, 'h21f8d, 'h10773, 'h10783, 'h10963, 'h10793, 'h10b63, 'h107a3, 'h10964, 'h107b3, 'h107c3, 'h10965, 'h107d3, 'h107e3, 'h10966, 'h107f3, 'h103bc, 'h10803, 'h10967, 'h10813, 'h21f8e, 'h21f8f, 'h21f8d, 'h10823, 'h10968, 'h10833, 'h10843, 'h10969, 'h10b63, 'h10853, 'h10863, 'h1096a, 'h10873, 'h10883, 'h1096b, 'h10893, 'h108a3, 'h1096c, 'h103bc, 'h108b3, 'h108c3, 'h1096d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d3, 'h106e3, 'h1096e, 'h10b73, 'h106f3, 'h10703, 'h1096f, 'h10713, 'h10723, 'h10970, 'h10733, 'h10743, 'h10971, 'h10753, 'h103bc, 'h10763, 'h10972, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10783, 'h10973, 'h10793, 'h10b73, 'h107a3, 'h10974, 'h107b3, 'h107c3, 'h10975, 'h107d3, 'h107e3, 'h10976, 'h107f3, 'h10803, 'h10977, 'h103bc, 'h10813, 'h10823, 'h10978, 'h21f8e, 'h21f8f, 'h21f8d, 'h10833, 'h10843, 'h10979, 'h10b73, 'h10853, 'h10863, 'h1097a, 'h10873, 'h10883, 'h1097b, 'h10893, 'h108a3, 'h1097c, 'h108b3, 'h103bc, 'h108c3, 'h1097d, 'h108d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1097e, 'h10b83, 'h106f3, 'h10703, 'h1097f, 'h10713, 'h10723, 'h10980, 'h10733, 'h10743, 'h10981, 'h10753, 'h10763, 'h10982, 'h103bc, 'h10773, 'h10783, 'h10983, 'h21f8e, 'h21f8f, 'h21f8d, 'h10793, 'h10b83, 'h107a3, 'h10984, 'h107b3, 'h107c3, 'h10985, 'h107d3, 'h107e3, 'h10986, 'h107f3, 'h10803, 'h10987, 'h10813, 'h103bc, 'h10823, 'h10988, 'h10833, 'h21f8e, 'h21f8f, 'h21f8d, 'h10843, 'h10989, 'h10b83, 'h10853, 'h10863, 'h1098a, 'h10873, 'h10883, 'h1098b, 'h10893, 'h108a3, 'h1098c, 'h108b3, 'h108c3, 'h1098d, 'h103bc, 'h108d3, 'h106e3, 'h1098e, 'h10b93, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f3, 'h10703, 'h1098f, 'h10713, 'h10723, 'h10990, 'h10733, 'h10743, 'h10991, 'h10753, 'h10763, 'h10992, 'h10773, 'h103bc, 'h10783, 'h10993, 'h10793, 'h10b93, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a3, 'h10994, 'h107b3, 'h107c3, 'h10995, 'h107d3, 'h107e3, 'h10996, 'h107f3, 'h10803, 'h10997, 'h10813, 'h10823, 'h10998, 'h103bc, 'h10833, 'h10843, 'h10999, 'h10b93, 'h21f8e, 'h21f8f, 'h21f8d, 'h10853, 'h10863, 'h1099a, 'h10873, 'h10883, 'h1099b, 'h10893, 'h108a3, 'h1099c, 'h108b3, 'h108c3, 'h1099d, 'h108d3, 'h103bc, 'h106e3, 'h1099e, 'h10ba3, 'h106f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10703, 'h1099f, 'h10713, 'h10723, 'h109a0, 'h10733, 'h10743, 'h109a1, 'h10753, 'h10763, 'h109a2, 'h10773, 'h10783, 'h109a3, 'h103bc, 'h10793, 'h10ba3, 'h107a3, 'h109a4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b3, 'h107c3, 'h109a5, 'h107d3, 'h107e3, 'h109a6, 'h107f3, 'h10803, 'h109a7, 'h10813, 'h10823, 'h109a8, 'h10833, 'h103bc, 'h10843, 'h109a9, 'h10ba3, 'h10853, 'h21f8e, 'h21f8f, 'h21f8d, 'h10863, 'h109aa, 'h10873, 'h10883, 'h109ab, 'h10893, 'h108a3, 'h109ac, 'h108b3, 'h108c3, 'h109ad, 'h108d3, 'h106e3, 'h109ae, 'h10bb3, 'h103bc, 'h106f3, 'h10703, 'h109af, 'h21f8e, 'h21f8f, 'h21f8d, 'h10713, 'h10723, 'h109b0, 'h10733, 'h10743, 'h109b1, 'h10753, 'h10763, 'h109b2, 'h10773, 'h10783, 'h109b3, 'h10793, 'h10bb3, 'h103bc, 'h107a3, 'h109b4, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c3, 'h109b5, 'h107d3, 'h107e3, 'h109b6, 'h107f3, 'h10803, 'h109b7, 'h10813, 'h10823, 'h109b8, 'h10833, 'h10843, 'h109b9, 'h10bb3, 'h103bc, 'h10853, 'h10863, 'h109ba, 'h21f8e, 'h21f8f, 'h21f8d, 'h10873, 'h10883, 'h109bb, 'h10893, 'h108a3, 'h109bc, 'h108b3, 'h108c3, 'h109bd, 'h108d3, 'h106e3, 'h109be, 'h10bc3, 'h106f3, 'h103bc, 'h10703, 'h109bf, 'h10713, 'h21f8e, 'h21f8f, 'h21f8d, 'h10723, 'h109c0, 'h10733, 'h10743, 'h109c1, 'h10753, 'h10763, 'h109c2, 'h10773, 'h10783, 'h109c3, 'h10793, 'h10bc3, 'h107a3, 'h109c4, 'h103bc, 'h107b3, 'h107c3, 'h109c5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d3, 'h107e3, 'h109c6, 'h107f3, 'h10803, 'h109c7, 'h10813, 'h10823, 'h109c8, 'h10833, 'h10843, 'h109c9, 'h10bc3, 'h10853, 'h103bc, 'h10863, 'h109ca, 'h10873, 'h21f8e, 'h21f8f, 'h21f8d, 'h10883, 'h109cb, 'h10893, 'h108a3, 'h109cc, 'h108b3, 'h108c3, 'h109cd, 'h108d3, 'h106e3, 'h109ce, 'h10bd3, 'h106f3, 'h10703, 'h109cf, 'h103bc, 'h10713, 'h10723, 'h109d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10733, 'h10743, 'h109d1, 'h10753, 'h10763, 'h109d2, 'h10773, 'h10783, 'h109d3, 'h10793, 'h10bd3, 'h107a3, 'h109d4, 'h107b3, 'h103bc, 'h107c3, 'h109d5, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e3, 'h109d6, 'h107f3, 'h10803, 'h109d7, 'h10813, 'h10823, 'h109d8, 'h10833, 'h10843, 'h109d9, 'h10bd3, 'h10853, 'h10863, 'h109da, 'h103bc, 'h10873, 'h10883, 'h109db, 'h21f8e, 'h21f8f, 'h21f8d, 'h10893, 'h108a3, 'h109dc, 'h108b3, 'h108c3, 'h109dd, 'h108d3, 'h106e3, 'h109de, 'h10be3, 'h106f3, 'h10703, 'h109df, 'h10713, 'h103bc, 'h10723, 'h109e0, 'h10733, 'h21f8e, 'h21f8f, 'h21f8d, 'h10743, 'h109e1, 'h10753, 'h10763, 'h109e2, 'h10773, 'h10783, 'h109e3, 'h10793, 'h10be3, 'h107a3, 'h109e4, 'h107b3, 'h107c3, 'h109e5, 'h103bc, 'h107d3, 'h107e3, 'h109e6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f3, 'h10803, 'h109e7, 'h10813, 'h10823, 'h109e8, 'h10833, 'h10843, 'h109e9, 'h10be3, 'h10853, 'h10863, 'h109ea, 'h10873, 'h103bc, 'h10883, 'h109eb, 'h10893, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a3, 'h109ec, 'h108b3, 'h108c3, 'h109ed, 'h108d3, 'h106e3, 'h109ee, 'h10bf3, 'h106f3, 'h10703, 'h109ef, 'h10713, 'h10723, 'h109f0, 'h103bc, 'h10733, 'h10743, 'h109f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10753, 'h10763, 'h109f2, 'h10773, 'h10783, 'h109f3, 'h10793, 'h10bf3, 'h107a3, 'h109f4, 'h107b3, 'h107c3, 'h109f5, 'h107d3, 'h103bc, 'h107e3, 'h109f6, 'h107f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10803, 'h109f7, 'h10813, 'h10823, 'h109f8, 'h10833, 'h10843, 'h109f9, 'h10bf3, 'h10853, 'h10863, 'h109fa, 'h10873, 'h10883, 'h109fb, 'h103bc, 'h10893, 'h108a3, 'h109fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b3, 'h108c3, 'h109fd, 'h108d3, 'h106e3, 'h109fe, 'h10c03, 'h106f3, 'h10703, 'h109ff, 'h10713, 'h10723, 'h10a00, 'h10733, 'h103bc, 'h10743, 'h10a01, 'h10753, 'h21f8e, 'h21f8f, 'h21f8d, 'h10763, 'h10a02, 'h10773, 'h10783, 'h10a03, 'h10793, 'h10c03, 'h107a3, 'h10a04, 'h107b3, 'h107c3, 'h10a05, 'h107d3, 'h107e3, 'h10a06, 'h103bc, 'h107f3, 'h10803, 'h10a07, 'h21f8e, 'h21f8f, 'h21f8d, 'h10813, 'h10823, 'h10a08, 'h10833, 'h10843, 'h10a09, 'h10c03, 'h10853, 'h10863, 'h10a0a, 'h10873, 'h10883, 'h10a0b, 'h10893, 'h103bc, 'h108a3, 'h10a0c, 'h108b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c3, 'h10a0d, 'h108d3, 'h106e3, 'h10a0e, 'h10c13, 'h106f3, 'h10703, 'h10a0f, 'h10713, 'h10723, 'h10a10, 'h10733, 'h10743, 'h10a11, 'h103bc, 'h10753, 'h10763, 'h10a12, 'h21f8e, 'h21f8f, 'h21f8d, 'h10773, 'h10783, 'h10a13, 'h10793, 'h10c13, 'h107a3, 'h10a14, 'h107b3, 'h107c3, 'h10a15, 'h107d3, 'h107e3, 'h10a16, 'h107f3, 'h103bc, 'h10803, 'h10a17, 'h10813, 'h21f8e, 'h21f8f, 'h21f8d, 'h10823, 'h10a18, 'h10833, 'h10843, 'h10a19, 'h10c13, 'h10853, 'h10863, 'h10a1a, 'h10873, 'h10883, 'h10a1b, 'h10893, 'h108a3, 'h10a1c, 'h103bc, 'h108b3, 'h108c3, 'h10a1d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d3, 'h106e3, 'h10a1e, 'h10c23, 'h106f3, 'h10703, 'h10a1f, 'h10713, 'h10723, 'h10a20, 'h10733, 'h10743, 'h10a21, 'h10753, 'h103bc, 'h10763, 'h10a22, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10783, 'h10a23, 'h10793, 'h10c23, 'h107a3, 'h10a24, 'h107b3, 'h107c3, 'h10a25, 'h107d3, 'h107e3, 'h10a26, 'h107f3, 'h10803, 'h10a27, 'h103bc, 'h10813, 'h10823, 'h10a28, 'h21f8e, 'h21f8f, 'h21f8d, 'h10833, 'h10843, 'h10a29, 'h10c23, 'h10853, 'h10863, 'h10a2a, 'h10873, 'h10883, 'h10a2b, 'h10893, 'h108a3, 'h10a2c, 'h108b3, 'h103bc, 'h108c3, 'h10a2d, 'h108d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h10a2e, 'h10c33, 'h106f3, 'h10703, 'h10a2f, 'h10713, 'h10723, 'h10a30, 'h10733, 'h10743, 'h10a31, 'h10753, 'h10763, 'h10a32, 'h103bc, 'h10773, 'h10783, 'h10a33, 'h21f8e, 'h21f8f, 'h21f8d, 'h10793, 'h10c33, 'h107a3, 'h10a34, 'h107b3, 'h107c3, 'h10a35, 'h107d3, 'h107e3, 'h10a36, 'h107f3, 'h10803, 'h10a37, 'h10813, 'h103bc, 'h10823, 'h10a38, 'h10833, 'h21f8e, 'h21f8f, 'h21f8d, 'h10843, 'h10a39, 'h10c33, 'h10853, 'h10863, 'h10a3a, 'h10873, 'h10883, 'h10a3b, 'h10893, 'h108a3, 'h10a3c, 'h108b3, 'h108c3, 'h10a3d, 'h103bc, 'h108d3, 'h106e3, 'h10a3e, 'h10c43, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f3, 'h10703, 'h10a3f, 'h10713, 'h10723, 'h10a40, 'h10733, 'h10743, 'h10a41, 'h10753, 'h10763, 'h10a42, 'h10773, 'h103bc, 'h10783, 'h10a43, 'h10793, 'h10c43, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a3, 'h10a44, 'h107b3, 'h107c3, 'h10a45, 'h107d3, 'h107e3, 'h10a46, 'h107f3, 'h10803, 'h10a47, 'h10813, 'h10823, 'h10a48, 'h103bc, 'h10833, 'h10843, 'h10a49, 'h10c43, 'h21f8e, 'h21f8f, 'h21f8d, 'h10853, 'h10863, 'h10a4a, 'h10873, 'h10883, 'h10a4b, 'h10893, 'h108a3, 'h10a4c, 'h108b3, 'h108c3, 'h10a4d, 'h108d3, 'h103bc, 'h106e3, 'h10a4e, 'h10c53, 'h106f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10703, 'h10a4f, 'h10713, 'h10723, 'h10a50, 'h10733, 'h10743, 'h10a51, 'h10753, 'h10763, 'h10a52, 'h10773, 'h10783, 'h10a53, 'h103bc, 'h10793, 'h10c53, 'h107a3, 'h10a54, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b3, 'h107c3, 'h10a55, 'h107d3, 'h107e3, 'h10a56, 'h107f3, 'h10803, 'h10a57, 'h10813, 'h10823, 'h10a58, 'h10833, 'h103bc, 'h10843, 'h10a59, 'h10c53, 'h10853, 'h21f8e, 'h21f8f, 'h21f8d, 'h10863, 'h10a5a, 'h10873, 'h10883, 'h10a5b, 'h10893, 'h108a3, 'h10a5c, 'h108b3, 'h108c3, 'h10a5d, 'h108d3, 'h106e3, 'h10a5e, 'h10c63, 'h103bc, 'h106f3, 'h10703, 'h10a5f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10713, 'h10723, 'h10a60, 'h10733, 'h10743, 'h10a61, 'h10753, 'h10763, 'h10a62, 'h10773, 'h10783, 'h10a63, 'h10793, 'h10c63, 'h103bc, 'h107a3, 'h10a64, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c3, 'h10a65, 'h107d3, 'h107e3, 'h10a66, 'h107f3, 'h10803, 'h10a67, 'h10813, 'h10823, 'h10a68, 'h10833, 'h10843, 'h10a69, 'h10c63, 'h103bc, 'h10853, 'h10863, 'h10a6a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10873, 'h10883, 'h10a6b, 'h10893, 'h108a3, 'h10a6c, 'h108b3, 'h108c3, 'h10a6d, 'h108d3, 'h106e3, 'h10a6e, 'h10c73, 'h106f3, 'h103bc, 'h10703, 'h10a6f, 'h10713, 'h21f8e, 'h21f8f, 'h21f8d, 'h10723, 'h10a70, 'h10733, 'h10743, 'h10a71, 'h10753, 'h10763, 'h10a72, 'h10773, 'h10783, 'h10a73, 'h10793, 'h10c73, 'h107a3, 'h10a74, 'h103bc, 'h107b3, 'h107c3, 'h10a75, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d3, 'h107e3, 'h10a76, 'h107f3, 'h10803, 'h10a77, 'h10813, 'h10823, 'h10a78, 'h10833, 'h10843, 'h10a79, 'h10c73, 'h10853, 'h103bc, 'h10863, 'h10a7a, 'h10873, 'h21f8e, 'h21f8f, 'h21f8d, 'h10883, 'h10a7b, 'h10893, 'h108a3, 'h10a7c, 'h108b3, 'h108c3, 'h10a7d, 'h108d3, 'h106e3, 'h10a7e, 'h10c83, 'h106f3, 'h10703, 'h10a7f, 'h103bc, 'h10713, 'h10723, 'h10a80, 'h21f8e, 'h21f8f, 'h21f8d, 'h10733, 'h10743, 'h10a81, 'h10753, 'h10763, 'h10a82, 'h10773, 'h10783, 'h10a83, 'h10793, 'h10c83, 'h107a3, 'h10a84, 'h107b3, 'h103bc, 'h107c3, 'h10a85, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e3, 'h10a86, 'h107f3, 'h10803, 'h10a87, 'h10813, 'h10823, 'h10a88, 'h10833, 'h10843, 'h10a89, 'h10c83, 'h10853, 'h10863, 'h10a8a, 'h103bc, 'h10873, 'h10883, 'h10a8b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10893, 'h108a3, 'h10a8c, 'h108b3, 'h108c3, 'h10a8d, 'h108d3, 'h106e3, 'h10a8e, 'h10c93, 'h106f3, 'h10703, 'h10a8f, 'h10713, 'h103bc, 'h10723, 'h10a90, 'h10733, 'h21f8e, 'h21f8f, 'h21f8d, 'h10743, 'h10a91, 'h10753, 'h10763, 'h10a92, 'h10773, 'h10783, 'h10a93, 'h10793, 'h10c93, 'h107a3, 'h10a94, 'h107b3, 'h107c3, 'h10a95, 'h103bc, 'h107d3, 'h107e3, 'h10a96, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f3, 'h10803, 'h10a97, 'h10813, 'h10823, 'h10a98, 'h10833, 'h10843, 'h10a99, 'h10c93, 'h10853, 'h10863, 'h10a9a, 'h10873, 'h103bc, 'h10883, 'h10a9b, 'h10893, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a3, 'h10a9c, 'h108b3, 'h108c3, 'h10a9d, 'h108d3, 'h106e3, 'h10a9e, 'h10ca3, 'h106f3, 'h10703, 'h10a9f, 'h10713, 'h10723, 'h10aa0, 'h103bc, 'h10733, 'h10743, 'h10aa1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10753, 'h10763, 'h10aa2, 'h10773, 'h10783, 'h10aa3, 'h10793, 'h10ca3, 'h107a3, 'h10aa4, 'h107b3, 'h107c3, 'h10aa5, 'h107d3, 'h103bc, 'h107e3, 'h10aa6, 'h107f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10803, 'h10aa7, 'h10813, 'h10823, 'h10aa8, 'h10833, 'h10843, 'h10aa9, 'h10ca3, 'h10853, 'h10863, 'h10aaa, 'h10873, 'h10883, 'h10aab, 'h103bc, 'h10893, 'h108a3, 'h10aac, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b3, 'h108c3, 'h10aad, 'h108d3, 'h106e3, 'h10aae, 'h10cb3, 'h106f3, 'h10703, 'h10aaf, 'h10713, 'h10723, 'h10ab0, 'h10733, 'h103bc, 'h10743, 'h10ab1, 'h10753, 'h21f8e, 'h21f8f, 'h21f8d, 'h10763, 'h10ab2, 'h10773, 'h10783, 'h10ab3, 'h10793, 'h10cb3, 'h107a3, 'h10ab4, 'h107b3, 'h107c3, 'h10ab5, 'h107d3, 'h107e3, 'h10ab6, 'h103bc, 'h107f3, 'h10803, 'h10ab7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10813, 'h10823, 'h10ab8, 'h10833, 'h10843, 'h10ab9, 'h10cb3, 'h10853, 'h10863, 'h10aba, 'h10873, 'h10883, 'h10abb, 'h10893, 'h103bc, 'h108a3, 'h10abc, 'h108b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c3, 'h10abd, 'h108d3, 'h106e3, 'h10abe, 'h10cc3, 'h106f3, 'h10703, 'h10abf, 'h10713, 'h10723, 'h10ac0, 'h10733, 'h10743, 'h10ac1, 'h103bc, 'h10753, 'h10763, 'h10ac2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10773, 'h10783, 'h10ac3, 'h10793, 'h10cc3, 'h107a3, 'h10ac4, 'h107b3, 'h107c3, 'h10ac5, 'h107d3, 'h107e3, 'h10ac6, 'h107f3, 'h103bc, 'h10803, 'h10ac7, 'h10813, 'h21f8e, 'h21f8f, 'h21f8d, 'h10823, 'h10ac8, 'h10833, 'h10843, 'h10ac9, 'h10cc3, 'h10853, 'h10863, 'h10aca, 'h10873, 'h10883, 'h10acb, 'h10893, 'h108a3, 'h10acc, 'h103bc, 'h108b3, 'h108c3, 'h10acd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d3, 'h106e3, 'h10ace, 'h10cd3, 'h106f3, 'h10703, 'h10acf, 'h10713, 'h10723, 'h10ad0, 'h10733, 'h10743, 'h10ad1, 'h10753, 'h103bc, 'h10763, 'h10ad2, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10783, 'h10ad3, 'h10793, 'h10cd3, 'h107a3, 'h10ad4, 'h107b3, 'h107c3, 'h10ad5, 'h107d3, 'h107e3, 'h10ad6, 'h107f3, 'h10803, 'h10ad7, 'h103bc, 'h10813, 'h10823, 'h10ad8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10833, 'h10843, 'h10ad9, 'h10cd3, 'h10853, 'h10863, 'h10ada, 'h10873, 'h10883, 'h10adb, 'h10893, 'h108a3, 'h10adc, 'h108b3, 'h103bc, 'h108c3, 'h10add, 'h108d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h108de, 'h10ae3, 'h106f3, 'h10703, 'h108df, 'h10713, 'h10723, 'h108e0, 'h10733, 'h10743, 'h108e1, 'h10753, 'h10763, 'h108e2, 'h103bc, 'h10773, 'h10783, 'h108e3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10793, 'h10ae3, 'h107a3, 'h108e4, 'h107b3, 'h107c3, 'h108e5, 'h107d3, 'h107e3, 'h108e6, 'h107f3, 'h10803, 'h108e7, 'h10813, 'h103bc, 'h10823, 'h108e8, 'h10833, 'h21f8e, 'h21f8f, 'h21f8d, 'h10843, 'h108e9, 'h10ae3, 'h10853, 'h10863, 'h108ea, 'h10873, 'h10883, 'h108eb, 'h10893, 'h108a3, 'h108ec, 'h108b3, 'h108c3, 'h108ed, 'h103bc, 'h108d3, 'h106e3, 'h108ee, 'h10af3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f3, 'h10703, 'h108ef, 'h10713, 'h10723, 'h108f0, 'h10733, 'h10743, 'h108f1, 'h10753, 'h10763, 'h108f2, 'h10773, 'h103bc, 'h10783, 'h108f3, 'h10793, 'h10af3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a3, 'h108f4, 'h107b3, 'h107c3, 'h108f5, 'h107d3, 'h107e3, 'h108f6, 'h107f3, 'h10803, 'h108f7, 'h10813, 'h10823, 'h108f8, 'h103bc, 'h10833, 'h10843, 'h108f9, 'h10af3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10853, 'h10863, 'h108fa, 'h10873, 'h10883, 'h108fb, 'h10893, 'h108a3, 'h108fc, 'h108b3, 'h108c3, 'h108fd, 'h108d3, 'h103bc, 'h106e3, 'h108fe, 'h10b03, 'h106f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10703, 'h108ff, 'h10713, 'h10723, 'h10900, 'h10733, 'h10743, 'h10901, 'h10753, 'h10763, 'h10902, 'h10773, 'h10783, 'h10903, 'h103bc, 'h10793, 'h10b03, 'h107a3, 'h10904, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b3, 'h107c3, 'h10905, 'h107d3, 'h107e3, 'h10906, 'h107f3, 'h10803, 'h10907, 'h10813, 'h10823, 'h10908, 'h10833, 'h103bc, 'h10843, 'h10909, 'h10b03, 'h10853, 'h21f8e, 'h21f8f, 'h21f8d, 'h10863, 'h1090a, 'h10873, 'h10883, 'h1090b, 'h10893, 'h108a3, 'h1090c, 'h108b3, 'h108c3, 'h1090d, 'h108d3, 'h106e3, 'h1090e, 'h10b13, 'h103bc, 'h106f3, 'h10703, 'h1090f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10713, 'h10723, 'h10910, 'h10733, 'h10743, 'h10911, 'h10753, 'h10763, 'h10912, 'h10773, 'h10783, 'h10913, 'h10793, 'h10b13, 'h103bc, 'h107a3, 'h10914, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c3, 'h10915, 'h107d3, 'h107e3, 'h10916, 'h107f3, 'h10803, 'h10917, 'h10813, 'h10823, 'h10918, 'h10833, 'h10843, 'h10919, 'h10b13, 'h103bc, 'h10853, 'h10863, 'h1091a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10873, 'h10883, 'h1091b, 'h10893, 'h108a3, 'h1091c, 'h108b3, 'h108c3, 'h1091d, 'h108d3, 'h106e3, 'h1091e, 'h10b23, 'h106f3, 'h103bc, 'h10703, 'h1091f, 'h10713, 'h21f8e, 'h21f8f, 'h21f8d, 'h10723, 'h10920, 'h10733, 'h10743, 'h10921, 'h10753, 'h10763, 'h10922, 'h10773, 'h10783, 'h10923, 'h10793, 'h10b23, 'h107a3, 'h10924, 'h103bc, 'h107b3, 'h107c3, 'h10925, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d3, 'h107e3, 'h10926, 'h107f3, 'h10803, 'h10927, 'h10813, 'h10823, 'h10928, 'h10833, 'h10843, 'h10929, 'h10b23, 'h10853, 'h103bc, 'h10863, 'h1092a, 'h10873, 'h21f8e, 'h21f8f, 'h21f8d, 'h10883, 'h1092b, 'h10893, 'h108a3, 'h1092c, 'h108b3, 'h108c3, 'h1092d, 'h108d3, 'h106e3, 'h1092e, 'h10b33, 'h106f3, 'h10703, 'h1092f, 'h103bc, 'h10713, 'h10723, 'h10930, 'h21f8e, 'h21f8f, 'h21f8d, 'h10733, 'h10743, 'h10931, 'h10753, 'h10763, 'h10932, 'h10773, 'h10783, 'h10933, 'h10793, 'h10b33, 'h107a3, 'h10934, 'h107b3, 'h103bc, 'h107c3, 'h10935, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e3, 'h10936, 'h107f3, 'h10803, 'h10937, 'h10813, 'h10823, 'h10938, 'h10833, 'h10843, 'h10939, 'h10b33, 'h10853, 'h10863, 'h1093a, 'h103bc, 'h10873, 'h10883, 'h1093b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10893, 'h108a3, 'h1093c, 'h108b3, 'h108c3, 'h1093d, 'h108d3, 'h106e3, 'h1093e, 'h10b43, 'h106f3, 'h10703, 'h1093f, 'h10713, 'h103bc, 'h10723, 'h10940, 'h10733, 'h21f8e, 'h21f8f, 'h21f8d, 'h10743, 'h10941, 'h10753, 'h10763, 'h10942, 'h10773, 'h10783, 'h10943, 'h10793, 'h10b43, 'h107a3, 'h10944, 'h107b3, 'h107c3, 'h10945, 'h103bc, 'h107d3, 'h107e3, 'h10946, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f3, 'h10803, 'h10947, 'h10813, 'h10823, 'h10948, 'h10833, 'h10843, 'h10949, 'h10b43, 'h10853, 'h10863, 'h1094a, 'h10873, 'h103bc, 'h10883, 'h1094b, 'h10893, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a3, 'h1094c, 'h108b3, 'h108c3, 'h1094d, 'h108d3, 'h106e3, 'h1094e, 'h10b53, 'h106f3, 'h10703, 'h1094f, 'h10713, 'h10723, 'h10950, 'h103bc, 'h10733, 'h10743, 'h10951, 'h21f8e, 'h21f8f, 'h21f8d, 'h10753, 'h10763, 'h10952, 'h10773, 'h10783, 'h10953, 'h10793, 'h10b53, 'h107a3, 'h10954, 'h107b3, 'h107c3, 'h10955, 'h107d3, 'h103bc, 'h107e3, 'h10956, 'h107f3, 'h21f8e, 'h21f8f};
	int DATA3 [3*SIZE-1:0] = {DATA2, DATA0};
	
endpackage
