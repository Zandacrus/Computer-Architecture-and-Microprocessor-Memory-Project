

package MATRIX_MULTIPLY_32_PKG_2;
	
	import MATRIX_MULTIPLY_32_PKG_1::DATA1;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h1072f, 'h1073f, 'h10a61, 'h1074f, 'h1075f, 'h10a62, 'h103bc, 'h1076f, 'h1077f, 'h10a63, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078f, 'h10c5f, 'h1079f, 'h10a64, 'h107af, 'h107bf, 'h10a65, 'h107cf, 'h107df, 'h10a66, 'h107ef, 'h107ff, 'h10a67, 'h1080f, 'h103bc, 'h1081f, 'h10a68, 'h1082f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083f, 'h10a69, 'h10c5f, 'h1084f, 'h1085f, 'h10a6a, 'h1086f, 'h1087f, 'h10a6b, 'h1088f, 'h1089f, 'h10a6c, 'h108af, 'h108bf, 'h10a6d, 'h103bc, 'h108cf, 'h106df, 'h10a6e, 'h10c6f, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ef, 'h106ff, 'h10a6f, 'h1070f, 'h1071f, 'h10a70, 'h1072f, 'h1073f, 'h10a71, 'h1074f, 'h1075f, 'h10a72, 'h1076f, 'h103bc, 'h1077f, 'h10a73, 'h1078f, 'h10c6f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079f, 'h10a74, 'h107af, 'h107bf, 'h10a75, 'h107cf, 'h107df, 'h10a76, 'h107ef, 'h107ff, 'h10a77, 'h1080f, 'h1081f, 'h10a78, 'h103bc, 'h1082f, 'h1083f, 'h10a79, 'h10c6f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084f, 'h1085f, 'h10a7a, 'h1086f, 'h1087f, 'h10a7b, 'h1088f, 'h1089f, 'h10a7c, 'h108af, 'h108bf, 'h10a7d, 'h108cf, 'h103bc, 'h106df, 'h10a7e, 'h10c7f, 'h106ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ff, 'h10a7f, 'h1070f, 'h1071f, 'h10a80, 'h1072f, 'h1073f, 'h10a81, 'h1074f, 'h1075f, 'h10a82, 'h1076f, 'h1077f, 'h10a83, 'h103bc, 'h1078f, 'h10c7f, 'h1079f, 'h10a84, 'h21f8e, 'h21f8f, 'h21f8d, 'h107af, 'h107bf, 'h10a85, 'h107cf, 'h107df, 'h10a86, 'h107ef, 'h107ff, 'h10a87, 'h1080f, 'h1081f, 'h10a88, 'h1082f, 'h103bc, 'h1083f, 'h10a89, 'h10c7f, 'h1084f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085f, 'h10a8a, 'h1086f, 'h1087f, 'h10a8b, 'h1088f, 'h1089f, 'h10a8c, 'h108af, 'h108bf, 'h10a8d, 'h108cf, 'h106df, 'h10a8e, 'h10c8f, 'h103bc, 'h106ef, 'h106ff, 'h10a8f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070f, 'h1071f, 'h10a90, 'h1072f, 'h1073f, 'h10a91, 'h1074f, 'h1075f, 'h10a92, 'h1076f, 'h1077f, 'h10a93, 'h1078f, 'h10c8f, 'h103bc, 'h1079f, 'h10a94, 'h107af, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bf, 'h10a95, 'h107cf, 'h107df, 'h10a96, 'h107ef, 'h107ff, 'h10a97, 'h1080f, 'h1081f, 'h10a98, 'h1082f, 'h1083f, 'h10a99, 'h10c8f, 'h103bc, 'h1084f, 'h1085f, 'h10a9a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086f, 'h1087f, 'h10a9b, 'h1088f, 'h1089f, 'h10a9c, 'h108af, 'h108bf, 'h10a9d, 'h108cf, 'h106df, 'h10a9e, 'h10c9f, 'h106ef, 'h103bc, 'h106ff, 'h10a9f, 'h1070f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071f, 'h10aa0, 'h1072f, 'h1073f, 'h10aa1, 'h1074f, 'h1075f, 'h10aa2, 'h1076f, 'h1077f, 'h10aa3, 'h1078f, 'h10c9f, 'h1079f, 'h10aa4, 'h103bc, 'h107af, 'h107bf, 'h10aa5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cf, 'h107df, 'h10aa6, 'h107ef, 'h107ff, 'h10aa7, 'h1080f, 'h1081f, 'h10aa8, 'h1082f, 'h1083f, 'h10aa9, 'h10c9f, 'h1084f, 'h103bc, 'h1085f, 'h10aaa, 'h1086f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087f, 'h10aab, 'h1088f, 'h1089f, 'h10aac, 'h108af, 'h108bf, 'h10aad, 'h108cf, 'h106df, 'h10aae, 'h10caf, 'h106ef, 'h106ff, 'h10aaf, 'h103bc, 'h1070f, 'h1071f, 'h10ab0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072f, 'h1073f, 'h10ab1, 'h1074f, 'h1075f, 'h10ab2, 'h1076f, 'h1077f, 'h10ab3, 'h1078f, 'h10caf, 'h1079f, 'h10ab4, 'h107af, 'h103bc, 'h107bf, 'h10ab5, 'h107cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h107df, 'h10ab6, 'h107ef, 'h107ff, 'h10ab7, 'h1080f, 'h1081f, 'h10ab8, 'h1082f, 'h1083f, 'h10ab9, 'h10caf, 'h1084f, 'h1085f, 'h10aba, 'h103bc, 'h1086f, 'h1087f, 'h10abb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088f, 'h1089f, 'h10abc, 'h108af, 'h108bf, 'h10abd, 'h108cf, 'h106df, 'h10abe, 'h10cbf, 'h106ef, 'h106ff, 'h10abf, 'h1070f, 'h103bc, 'h1071f, 'h10ac0, 'h1072f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073f, 'h10ac1, 'h1074f, 'h1075f, 'h10ac2, 'h1076f, 'h1077f, 'h10ac3, 'h1078f, 'h10cbf, 'h1079f, 'h10ac4, 'h107af, 'h107bf, 'h10ac5, 'h103bc, 'h107cf, 'h107df, 'h10ac6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ef, 'h107ff, 'h10ac7, 'h1080f, 'h1081f, 'h10ac8, 'h1082f, 'h1083f, 'h10ac9, 'h10cbf, 'h1084f, 'h1085f, 'h10aca, 'h1086f, 'h103bc, 'h1087f, 'h10acb, 'h1088f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089f, 'h10acc, 'h108af, 'h108bf, 'h10acd, 'h108cf, 'h106df, 'h10ace, 'h10ccf, 'h106ef, 'h106ff, 'h10acf, 'h1070f, 'h1071f, 'h10ad0, 'h103bc, 'h1072f, 'h1073f, 'h10ad1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074f, 'h1075f, 'h10ad2, 'h1076f, 'h1077f, 'h10ad3, 'h1078f, 'h10ccf, 'h1079f, 'h10ad4, 'h107af, 'h107bf, 'h10ad5, 'h107cf, 'h103bc, 'h107df, 'h10ad6, 'h107ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ff, 'h10ad7, 'h1080f, 'h1081f, 'h10ad8, 'h1082f, 'h1083f, 'h10ad9, 'h10ccf, 'h1084f, 'h1085f, 'h10ada, 'h1086f, 'h1087f, 'h10adb, 'h103bc, 'h1088f, 'h1089f, 'h10adc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108af, 'h108bf, 'h10add, 'h108cf, 'h106df, 'h108de, 'h10adf, 'h106ef, 'h106ff, 'h108df, 'h1070f, 'h1071f, 'h108e0, 'h1072f, 'h103bc, 'h1073f, 'h108e1, 'h1074f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075f, 'h108e2, 'h1076f, 'h1077f, 'h108e3, 'h1078f, 'h10adf, 'h1079f, 'h108e4, 'h107af, 'h107bf, 'h108e5, 'h107cf, 'h107df, 'h108e6, 'h103bc, 'h107ef, 'h107ff, 'h108e7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080f, 'h1081f, 'h108e8, 'h1082f, 'h1083f, 'h108e9, 'h10adf, 'h1084f, 'h1085f, 'h108ea, 'h1086f, 'h1087f, 'h108eb, 'h1088f, 'h103bc, 'h1089f, 'h108ec, 'h108af, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bf, 'h108ed, 'h108cf, 'h106df, 'h108ee, 'h10aef, 'h106ef, 'h106ff, 'h108ef, 'h1070f, 'h1071f, 'h108f0, 'h1072f, 'h1073f, 'h108f1, 'h103bc, 'h1074f, 'h1075f, 'h108f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076f, 'h1077f, 'h108f3, 'h1078f, 'h10aef, 'h1079f, 'h108f4, 'h107af, 'h107bf, 'h108f5, 'h107cf, 'h107df, 'h108f6, 'h107ef, 'h103bc, 'h107ff, 'h108f7, 'h1080f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081f, 'h108f8, 'h1082f, 'h1083f, 'h108f9, 'h10aef, 'h1084f, 'h1085f, 'h108fa, 'h1086f, 'h1087f, 'h108fb, 'h1088f, 'h1089f, 'h108fc, 'h103bc, 'h108af, 'h108bf, 'h108fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cf, 'h106df, 'h108fe, 'h10aff, 'h106ef, 'h106ff, 'h108ff, 'h1070f, 'h1071f, 'h10900, 'h1072f, 'h1073f, 'h10901, 'h1074f, 'h103bc, 'h1075f, 'h10902, 'h1076f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077f, 'h10903, 'h1078f, 'h10aff, 'h1079f, 'h10904, 'h107af, 'h107bf, 'h10905, 'h107cf, 'h107df, 'h10906, 'h107ef, 'h107ff, 'h10907, 'h103bc, 'h1080f, 'h1081f, 'h10908, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082f, 'h1083f, 'h10909, 'h10aff, 'h1084f, 'h1085f, 'h1090a, 'h1086f, 'h1087f, 'h1090b, 'h1088f, 'h1089f, 'h1090c, 'h108af, 'h103bc, 'h108bf, 'h1090d, 'h108cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1090e, 'h10b0f, 'h106ef, 'h106ff, 'h1090f, 'h1070f, 'h1071f, 'h10910, 'h1072f, 'h1073f, 'h10911, 'h1074f, 'h1075f, 'h10912, 'h103bc, 'h1076f, 'h1077f, 'h10913, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078f, 'h10b0f, 'h1079f, 'h10914, 'h107af, 'h107bf, 'h10915, 'h107cf, 'h107df, 'h10916, 'h107ef, 'h107ff, 'h10917, 'h1080f, 'h103bc, 'h1081f, 'h10918, 'h1082f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083f, 'h10919, 'h10b0f, 'h1084f, 'h1085f, 'h1091a, 'h1086f, 'h1087f, 'h1091b, 'h1088f, 'h1089f, 'h1091c, 'h108af, 'h108bf, 'h1091d, 'h103bc, 'h108cf, 'h106df, 'h1091e, 'h10b1f, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ef, 'h106ff, 'h1091f, 'h1070f, 'h1071f, 'h10920, 'h1072f, 'h1073f, 'h10921, 'h1074f, 'h1075f, 'h10922, 'h1076f, 'h103bc, 'h1077f, 'h10923, 'h1078f, 'h10b1f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079f, 'h10924, 'h107af, 'h107bf, 'h10925, 'h107cf, 'h107df, 'h10926, 'h107ef, 'h107ff, 'h10927, 'h1080f, 'h1081f, 'h10928, 'h103bc, 'h1082f, 'h1083f, 'h10929, 'h10b1f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084f, 'h1085f, 'h1092a, 'h1086f, 'h1087f, 'h1092b, 'h1088f, 'h1089f, 'h1092c, 'h108af, 'h108bf, 'h1092d, 'h108cf, 'h103bc, 'h106df, 'h1092e, 'h10b2f, 'h106ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ff, 'h1092f, 'h1070f, 'h1071f, 'h10930, 'h1072f, 'h1073f, 'h10931, 'h1074f, 'h1075f, 'h10932, 'h1076f, 'h1077f, 'h10933, 'h103bc, 'h1078f, 'h10b2f, 'h1079f, 'h10934, 'h21f8e, 'h21f8f, 'h21f8d, 'h107af, 'h107bf, 'h10935, 'h107cf, 'h107df, 'h10936, 'h107ef, 'h107ff, 'h10937, 'h1080f, 'h1081f, 'h10938, 'h1082f, 'h103bc, 'h1083f, 'h10939, 'h10b2f, 'h1084f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085f, 'h1093a, 'h1086f, 'h1087f, 'h1093b, 'h1088f, 'h1089f, 'h1093c, 'h108af, 'h108bf, 'h1093d, 'h108cf, 'h106df, 'h1093e, 'h10b3f, 'h103bc, 'h106ef, 'h106ff, 'h1093f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070f, 'h1071f, 'h10940, 'h1072f, 'h1073f, 'h10941, 'h1074f, 'h1075f, 'h10942, 'h1076f, 'h1077f, 'h10943, 'h1078f, 'h10b3f, 'h103bc, 'h1079f, 'h10944, 'h107af, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bf, 'h10945, 'h107cf, 'h107df, 'h10946, 'h107ef, 'h107ff, 'h10947, 'h1080f, 'h1081f, 'h10948, 'h1082f, 'h1083f, 'h10949, 'h10b3f, 'h103bc, 'h1084f, 'h1085f, 'h1094a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086f, 'h1087f, 'h1094b, 'h1088f, 'h1089f, 'h1094c, 'h108af, 'h108bf, 'h1094d, 'h108cf, 'h106df, 'h1094e, 'h10b4f, 'h106ef, 'h103bc, 'h106ff, 'h1094f, 'h1070f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071f, 'h10950, 'h1072f, 'h1073f, 'h10951, 'h1074f, 'h1075f, 'h10952, 'h1076f, 'h1077f, 'h10953, 'h1078f, 'h10b4f, 'h1079f, 'h10954, 'h103bc, 'h107af, 'h107bf, 'h10955, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cf, 'h107df, 'h10956, 'h107ef, 'h107ff, 'h10957, 'h1080f, 'h1081f, 'h10958, 'h1082f, 'h1083f, 'h10959, 'h10b4f, 'h1084f, 'h103bc, 'h1085f, 'h1095a, 'h1086f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087f, 'h1095b, 'h1088f, 'h1089f, 'h1095c, 'h108af, 'h108bf, 'h1095d, 'h108cf, 'h106df, 'h1095e, 'h10b5f, 'h106ef, 'h106ff, 'h1095f, 'h103bc, 'h1070f, 'h1071f, 'h10960, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072f, 'h1073f, 'h10961, 'h1074f, 'h1075f, 'h10962, 'h1076f, 'h1077f, 'h10963, 'h1078f, 'h10b5f, 'h1079f, 'h10964, 'h107af, 'h103bc, 'h107bf, 'h10965, 'h107cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h107df, 'h10966, 'h107ef, 'h107ff, 'h10967, 'h1080f, 'h1081f, 'h10968, 'h1082f, 'h1083f, 'h10969, 'h10b5f, 'h1084f, 'h1085f, 'h1096a, 'h103bc, 'h1086f, 'h1087f, 'h1096b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088f, 'h1089f, 'h1096c, 'h108af, 'h108bf, 'h1096d, 'h108cf, 'h106df, 'h1096e, 'h10b6f, 'h106ef, 'h106ff, 'h1096f, 'h1070f, 'h103bc, 'h1071f, 'h10970, 'h1072f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073f, 'h10971, 'h1074f, 'h1075f, 'h10972, 'h1076f, 'h1077f, 'h10973, 'h1078f, 'h10b6f, 'h1079f, 'h10974, 'h107af, 'h107bf, 'h10975, 'h103bc, 'h107cf, 'h107df, 'h10976, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ef, 'h107ff, 'h10977, 'h1080f, 'h1081f, 'h10978, 'h1082f, 'h1083f, 'h10979, 'h10b6f, 'h1084f, 'h1085f, 'h1097a, 'h1086f, 'h103bc, 'h1087f, 'h1097b, 'h1088f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089f, 'h1097c, 'h108af, 'h108bf, 'h1097d, 'h108cf, 'h106df, 'h1097e, 'h10b7f, 'h106ef, 'h106ff, 'h1097f, 'h1070f, 'h1071f, 'h10980, 'h103bc, 'h1072f, 'h1073f, 'h10981, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074f, 'h1075f, 'h10982, 'h1076f, 'h1077f, 'h10983, 'h1078f, 'h10b7f, 'h1079f, 'h10984, 'h107af, 'h107bf, 'h10985, 'h107cf, 'h103bc, 'h107df, 'h10986, 'h107ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ff, 'h10987, 'h1080f, 'h1081f, 'h10988, 'h1082f, 'h1083f, 'h10989, 'h10b7f, 'h1084f, 'h1085f, 'h1098a, 'h1086f, 'h1087f, 'h1098b, 'h103bc, 'h1088f, 'h1089f, 'h1098c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108af, 'h108bf, 'h1098d, 'h108cf, 'h106df, 'h1098e, 'h10b8f, 'h106ef, 'h106ff, 'h1098f, 'h1070f, 'h1071f, 'h10990, 'h1072f, 'h103bc, 'h1073f, 'h10991, 'h1074f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075f, 'h10992, 'h1076f, 'h1077f, 'h10993, 'h1078f, 'h10b8f, 'h1079f, 'h10994, 'h107af, 'h107bf, 'h10995, 'h107cf, 'h107df, 'h10996, 'h103bc, 'h107ef, 'h107ff, 'h10997, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080f, 'h1081f, 'h10998, 'h1082f, 'h1083f, 'h10999, 'h10b8f, 'h1084f, 'h1085f, 'h1099a, 'h1086f, 'h1087f, 'h1099b, 'h1088f, 'h103bc, 'h1089f, 'h1099c, 'h108af, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bf, 'h1099d, 'h108cf, 'h106df, 'h1099e, 'h10b9f, 'h106ef, 'h106ff, 'h1099f, 'h1070f, 'h1071f, 'h109a0, 'h1072f, 'h1073f, 'h109a1, 'h103bc, 'h1074f, 'h1075f, 'h109a2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076f, 'h1077f, 'h109a3, 'h1078f, 'h10b9f, 'h1079f, 'h109a4, 'h107af, 'h107bf, 'h109a5, 'h107cf, 'h107df, 'h109a6, 'h107ef, 'h103bc, 'h107ff, 'h109a7, 'h1080f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081f, 'h109a8, 'h1082f, 'h1083f, 'h109a9, 'h10b9f, 'h1084f, 'h1085f, 'h109aa, 'h1086f, 'h1087f, 'h109ab, 'h1088f, 'h1089f, 'h109ac, 'h103bc, 'h108af, 'h108bf, 'h109ad, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cf, 'h106df, 'h109ae, 'h10baf, 'h106ef, 'h106ff, 'h109af, 'h1070f, 'h1071f, 'h109b0, 'h1072f, 'h1073f, 'h109b1, 'h1074f, 'h103bc, 'h1075f, 'h109b2, 'h1076f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077f, 'h109b3, 'h1078f, 'h10baf, 'h1079f, 'h109b4, 'h107af, 'h107bf, 'h109b5, 'h107cf, 'h107df, 'h109b6, 'h107ef, 'h107ff, 'h109b7, 'h103bc, 'h1080f, 'h1081f, 'h109b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082f, 'h1083f, 'h109b9, 'h10baf, 'h1084f, 'h1085f, 'h109ba, 'h1086f, 'h1087f, 'h109bb, 'h1088f, 'h1089f, 'h109bc, 'h108af, 'h103bc, 'h108bf, 'h109bd, 'h108cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h109be, 'h10bbf, 'h106ef, 'h106ff, 'h109bf, 'h1070f, 'h1071f, 'h109c0, 'h1072f, 'h1073f, 'h109c1, 'h1074f, 'h1075f, 'h109c2, 'h103bc, 'h1076f, 'h1077f, 'h109c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078f, 'h10bbf, 'h1079f, 'h109c4, 'h107af, 'h107bf, 'h109c5, 'h107cf, 'h107df, 'h109c6, 'h107ef, 'h107ff, 'h109c7, 'h1080f, 'h103bc, 'h1081f, 'h109c8, 'h1082f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083f, 'h109c9, 'h10bbf, 'h1084f, 'h1085f, 'h109ca, 'h1086f, 'h1087f, 'h109cb, 'h1088f, 'h1089f, 'h109cc, 'h108af, 'h108bf, 'h109cd, 'h103bc, 'h108cf, 'h106df, 'h109ce, 'h10bcf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ef, 'h106ff, 'h109cf, 'h1070f, 'h1071f, 'h109d0, 'h1072f, 'h1073f, 'h109d1, 'h1074f, 'h1075f, 'h109d2, 'h1076f, 'h103bc, 'h1077f, 'h109d3, 'h1078f, 'h10bcf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079f, 'h109d4, 'h107af, 'h107bf, 'h109d5, 'h107cf, 'h107df, 'h109d6, 'h107ef, 'h107ff, 'h109d7, 'h1080f, 'h1081f, 'h109d8, 'h103bc, 'h1082f, 'h1083f, 'h109d9, 'h10bcf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084f, 'h1085f, 'h109da, 'h1086f, 'h1087f, 'h109db, 'h1088f, 'h1089f, 'h109dc, 'h108af, 'h108bf, 'h109dd, 'h108cf, 'h103bc, 'h106df, 'h109de, 'h10bdf, 'h106ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ff, 'h109df, 'h1070f, 'h1071f, 'h109e0, 'h1072f, 'h1073f, 'h109e1, 'h1074f, 'h1075f, 'h109e2, 'h1076f, 'h1077f, 'h109e3, 'h103bc, 'h1078f, 'h10bdf, 'h1079f, 'h109e4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107af, 'h107bf, 'h109e5, 'h107cf, 'h107df, 'h109e6, 'h107ef, 'h107ff, 'h109e7, 'h1080f, 'h1081f, 'h109e8, 'h1082f, 'h103bc, 'h1083f, 'h109e9, 'h10bdf, 'h1084f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085f, 'h109ea, 'h1086f, 'h1087f, 'h109eb, 'h1088f, 'h1089f, 'h109ec, 'h108af, 'h108bf, 'h109ed, 'h108cf, 'h106df, 'h109ee, 'h10bef, 'h103bc, 'h106ef, 'h106ff, 'h109ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070f, 'h1071f, 'h109f0, 'h1072f, 'h1073f, 'h109f1, 'h1074f, 'h1075f, 'h109f2, 'h1076f, 'h1077f, 'h109f3, 'h1078f, 'h10bef, 'h103bc, 'h1079f, 'h109f4, 'h107af, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bf, 'h109f5, 'h107cf, 'h107df, 'h109f6, 'h107ef, 'h107ff, 'h109f7, 'h1080f, 'h1081f, 'h109f8, 'h1082f, 'h1083f, 'h109f9, 'h10bef, 'h103bc, 'h1084f, 'h1085f, 'h109fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086f, 'h1087f, 'h109fb, 'h1088f, 'h1089f, 'h109fc, 'h108af, 'h108bf, 'h109fd, 'h108cf, 'h106df, 'h109fe, 'h10bff, 'h106ef, 'h103bc, 'h106ff, 'h109ff, 'h1070f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071f, 'h10a00, 'h1072f, 'h1073f, 'h10a01, 'h1074f, 'h1075f, 'h10a02, 'h1076f, 'h1077f, 'h10a03, 'h1078f, 'h10bff, 'h1079f, 'h10a04, 'h103bc, 'h107af, 'h107bf, 'h10a05, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cf, 'h107df, 'h10a06, 'h107ef, 'h107ff, 'h10a07, 'h1080f, 'h1081f, 'h10a08, 'h1082f, 'h1083f, 'h10a09, 'h10bff, 'h1084f, 'h103bc, 'h1085f, 'h10a0a, 'h1086f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087f, 'h10a0b, 'h1088f, 'h1089f, 'h10a0c, 'h108af, 'h108bf, 'h10a0d, 'h108cf, 'h106df, 'h10a0e, 'h10c0f, 'h106ef, 'h106ff, 'h10a0f, 'h103bc, 'h1070f, 'h1071f, 'h10a10, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072f, 'h1073f, 'h10a11, 'h1074f, 'h1075f, 'h10a12, 'h1076f, 'h1077f, 'h10a13, 'h1078f, 'h10c0f, 'h1079f, 'h10a14, 'h107af, 'h103bc, 'h107bf, 'h10a15, 'h107cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h107df, 'h10a16, 'h107ef, 'h107ff, 'h10a17, 'h1080f, 'h1081f, 'h10a18, 'h1082f, 'h1083f, 'h10a19, 'h10c0f, 'h1084f, 'h1085f, 'h10a1a, 'h103bc, 'h1086f, 'h1087f, 'h10a1b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088f, 'h1089f, 'h10a1c, 'h108af, 'h108bf, 'h10a1d, 'h108cf, 'h106df, 'h10a1e, 'h10c1f, 'h106ef, 'h106ff, 'h10a1f, 'h1070f, 'h103bc, 'h1071f, 'h10a20, 'h1072f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073f, 'h10a21, 'h1074f, 'h1075f, 'h10a22, 'h1076f, 'h1077f, 'h10a23, 'h1078f, 'h10c1f, 'h1079f, 'h10a24, 'h107af, 'h107bf, 'h10a25, 'h103bc, 'h107cf, 'h107df, 'h10a26, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ef, 'h107ff, 'h10a27, 'h1080f, 'h1081f, 'h10a28, 'h1082f, 'h1083f, 'h10a29, 'h10c1f, 'h1084f, 'h1085f, 'h10a2a, 'h1086f, 'h103bc, 'h1087f, 'h10a2b, 'h1088f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089f, 'h10a2c, 'h108af, 'h108bf, 'h10a2d, 'h108cf, 'h106df, 'h10a2e, 'h10c2f, 'h106ef, 'h106ff, 'h10a2f, 'h1070f, 'h1071f, 'h10a30, 'h103bc, 'h1072f, 'h1073f, 'h10a31, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074f, 'h1075f, 'h10a32, 'h1076f, 'h1077f, 'h10a33, 'h1078f, 'h10c2f, 'h1079f, 'h10a34, 'h107af, 'h107bf, 'h10a35, 'h107cf, 'h103bc, 'h107df, 'h10a36, 'h107ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ff, 'h10a37, 'h1080f, 'h1081f, 'h10a38, 'h1082f, 'h1083f, 'h10a39, 'h10c2f, 'h1084f, 'h1085f, 'h10a3a, 'h1086f, 'h1087f, 'h10a3b, 'h103bc, 'h1088f, 'h1089f, 'h10a3c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108af, 'h108bf, 'h10a3d, 'h108cf, 'h106df, 'h10a3e, 'h10c3f, 'h106ef, 'h106ff, 'h10a3f, 'h1070f, 'h1071f, 'h10a40, 'h1072f, 'h103bc, 'h1073f, 'h10a41, 'h1074f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075f, 'h10a42, 'h1076f, 'h1077f, 'h10a43, 'h1078f, 'h10c3f, 'h1079f, 'h10a44, 'h107af, 'h107bf, 'h10a45, 'h107cf, 'h107df, 'h10a46, 'h103bc, 'h107ef, 'h107ff, 'h10a47, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080f, 'h1081f, 'h10a48, 'h1082f, 'h1083f, 'h10a49, 'h10c3f, 'h1084f, 'h1085f, 'h10a4a, 'h1086f, 'h1087f, 'h10a4b, 'h1088f, 'h103bc, 'h1089f, 'h10a4c, 'h108af, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bf, 'h10a4d, 'h108cf, 'h106df, 'h10a4e, 'h10c4f, 'h106ef, 'h106ff, 'h10a4f, 'h1070f, 'h1071f, 'h10a50, 'h1072f, 'h1073f, 'h10a51, 'h103bc, 'h1074f, 'h1075f, 'h10a52, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076f, 'h1077f, 'h10a53, 'h1078f, 'h10c4f, 'h1079f, 'h10a54, 'h107af, 'h107bf, 'h10a55, 'h107cf, 'h107df, 'h10a56, 'h107ef, 'h103bc, 'h107ff, 'h10a57, 'h1080f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081f, 'h10a58, 'h1082f, 'h1083f, 'h10a59, 'h10c4f, 'h1084f, 'h1085f, 'h10a5a, 'h1086f, 'h1087f, 'h10a5b, 'h1088f, 'h1089f, 'h10a5c, 'h103bc, 'h108af, 'h108bf, 'h10a5d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cf, 'h106df, 'h10a5e, 'h10c5f, 'h106ef, 'h106ff, 'h10a5f, 'h1070f, 'h1071f, 'h10a60, 'h1072f, 'h1073f, 'h10a61, 'h1074f, 'h103bc, 'h1075f, 'h10a62, 'h1076f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077f, 'h10a63, 'h1078f, 'h10c5f, 'h1079f, 'h10a64, 'h107af, 'h107bf, 'h10a65, 'h107cf, 'h107df, 'h10a66, 'h107ef, 'h107ff, 'h10a67, 'h103bc, 'h1080f, 'h1081f, 'h10a68, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082f, 'h1083f, 'h10a69, 'h10c5f, 'h1084f, 'h1085f, 'h10a6a, 'h1086f, 'h1087f, 'h10a6b, 'h1088f, 'h1089f, 'h10a6c, 'h108af, 'h103bc, 'h108bf, 'h10a6d, 'h108cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h10a6e, 'h10c6f, 'h106ef, 'h106ff, 'h10a6f, 'h1070f, 'h1071f, 'h10a70, 'h1072f, 'h1073f, 'h10a71, 'h1074f, 'h1075f, 'h10a72, 'h103bc, 'h1076f, 'h1077f, 'h10a73, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078f, 'h10c6f, 'h1079f, 'h10a74, 'h107af, 'h107bf, 'h10a75, 'h107cf, 'h107df, 'h10a76, 'h107ef, 'h107ff, 'h10a77, 'h1080f, 'h103bc, 'h1081f, 'h10a78, 'h1082f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083f, 'h10a79, 'h10c6f, 'h1084f, 'h1085f, 'h10a7a, 'h1086f, 'h1087f, 'h10a7b, 'h1088f, 'h1089f, 'h10a7c, 'h108af, 'h108bf, 'h10a7d, 'h103bc, 'h108cf, 'h106df, 'h10a7e, 'h10c7f, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ef, 'h106ff, 'h10a7f, 'h1070f, 'h1071f, 'h10a80, 'h1072f, 'h1073f, 'h10a81, 'h1074f, 'h1075f, 'h10a82, 'h1076f, 'h103bc, 'h1077f, 'h10a83, 'h1078f, 'h10c7f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079f, 'h10a84, 'h107af, 'h107bf, 'h10a85, 'h107cf, 'h107df, 'h10a86, 'h107ef, 'h107ff, 'h10a87, 'h1080f, 'h1081f, 'h10a88, 'h103bc, 'h1082f, 'h1083f, 'h10a89, 'h10c7f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084f, 'h1085f, 'h10a8a, 'h1086f, 'h1087f, 'h10a8b, 'h1088f, 'h1089f, 'h10a8c, 'h108af, 'h108bf, 'h10a8d, 'h108cf, 'h103bc, 'h106df, 'h10a8e, 'h10c8f, 'h106ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ff, 'h10a8f, 'h1070f, 'h1071f, 'h10a90, 'h1072f, 'h1073f, 'h10a91, 'h1074f, 'h1075f, 'h10a92, 'h1076f, 'h1077f, 'h10a93, 'h103bc, 'h1078f, 'h10c8f, 'h1079f, 'h10a94, 'h21f8e, 'h21f8f, 'h21f8d, 'h107af, 'h107bf, 'h10a95, 'h107cf, 'h107df, 'h10a96, 'h107ef, 'h107ff, 'h10a97, 'h1080f, 'h1081f, 'h10a98, 'h1082f, 'h103bc, 'h1083f, 'h10a99, 'h10c8f, 'h1084f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085f, 'h10a9a, 'h1086f, 'h1087f, 'h10a9b, 'h1088f, 'h1089f, 'h10a9c, 'h108af, 'h108bf, 'h10a9d, 'h108cf, 'h106df, 'h10a9e, 'h10c9f, 'h103bc, 'h106ef, 'h106ff, 'h10a9f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070f, 'h1071f, 'h10aa0, 'h1072f, 'h1073f, 'h10aa1, 'h1074f, 'h1075f, 'h10aa2, 'h1076f, 'h1077f, 'h10aa3, 'h1078f, 'h10c9f, 'h103bc, 'h1079f, 'h10aa4, 'h107af, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bf, 'h10aa5, 'h107cf, 'h107df, 'h10aa6, 'h107ef, 'h107ff, 'h10aa7, 'h1080f, 'h1081f, 'h10aa8, 'h1082f, 'h1083f, 'h10aa9, 'h10c9f, 'h103bc, 'h1084f, 'h1085f, 'h10aaa, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086f, 'h1087f, 'h10aab, 'h1088f, 'h1089f, 'h10aac, 'h108af, 'h108bf, 'h10aad, 'h108cf, 'h106df, 'h10aae, 'h10caf, 'h106ef, 'h103bc, 'h106ff, 'h10aaf, 'h1070f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071f, 'h10ab0, 'h1072f, 'h1073f, 'h10ab1, 'h1074f, 'h1075f, 'h10ab2, 'h1076f, 'h1077f, 'h10ab3, 'h1078f, 'h10caf, 'h1079f, 'h10ab4, 'h103bc, 'h107af, 'h107bf, 'h10ab5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cf, 'h107df, 'h10ab6, 'h107ef, 'h107ff, 'h10ab7, 'h1080f, 'h1081f, 'h10ab8, 'h1082f, 'h1083f, 'h10ab9, 'h10caf, 'h1084f, 'h103bc, 'h1085f, 'h10aba, 'h1086f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087f, 'h10abb, 'h1088f, 'h1089f, 'h10abc, 'h108af, 'h108bf, 'h10abd, 'h108cf, 'h106df, 'h10abe, 'h10cbf, 'h106ef, 'h106ff, 'h10abf, 'h103bc, 'h1070f, 'h1071f, 'h10ac0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072f, 'h1073f, 'h10ac1, 'h1074f, 'h1075f, 'h10ac2, 'h1076f, 'h1077f, 'h10ac3, 'h1078f, 'h10cbf, 'h1079f, 'h10ac4, 'h107af, 'h103bc, 'h107bf, 'h10ac5, 'h107cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h107df, 'h10ac6, 'h107ef, 'h107ff, 'h10ac7, 'h1080f, 'h1081f, 'h10ac8, 'h1082f, 'h1083f, 'h10ac9, 'h10cbf, 'h1084f, 'h1085f, 'h10aca, 'h103bc, 'h1086f, 'h1087f, 'h10acb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088f, 'h1089f, 'h10acc, 'h108af, 'h108bf, 'h10acd, 'h108cf, 'h106df, 'h10ace, 'h10ccf, 'h106ef, 'h106ff, 'h10acf, 'h1070f, 'h103bc, 'h1071f, 'h10ad0, 'h1072f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073f, 'h10ad1, 'h1074f, 'h1075f, 'h10ad2, 'h1076f, 'h1077f, 'h10ad3, 'h1078f, 'h10ccf, 'h1079f, 'h10ad4, 'h107af, 'h107bf, 'h10ad5, 'h103bc, 'h107cf, 'h107df, 'h10ad6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ef, 'h107ff, 'h10ad7, 'h1080f, 'h1081f, 'h10ad8, 'h1082f, 'h1083f, 'h10ad9, 'h10ccf, 'h1084f, 'h1085f, 'h10ada, 'h1086f, 'h103bc, 'h1087f, 'h10adb, 'h1088f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089f, 'h10adc, 'h108af, 'h108bf, 'h10add, 'h108cf, 'h106e0, 'h108de, 'h10ae0, 'h106f0, 'h10700, 'h108df, 'h10710, 'h10720, 'h108e0, 'h103bc, 'h10730, 'h10740, 'h108e1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10750, 'h10760, 'h108e2, 'h10770, 'h10780, 'h108e3, 'h10790, 'h10ae0, 'h107a0, 'h108e4, 'h107b0, 'h107c0, 'h108e5, 'h107d0, 'h103bc, 'h107e0, 'h108e6, 'h107f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10800, 'h108e7, 'h10810, 'h10820, 'h108e8, 'h10830, 'h10840, 'h108e9, 'h10ae0, 'h10850, 'h10860, 'h108ea, 'h10870, 'h10880, 'h108eb, 'h103bc, 'h10890, 'h108a0, 'h108ec, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b0, 'h108c0, 'h108ed, 'h108d0, 'h106e0, 'h108ee, 'h10af0, 'h106f0, 'h10700, 'h108ef, 'h10710, 'h10720, 'h108f0, 'h10730, 'h103bc, 'h10740, 'h108f1, 'h10750, 'h21f8e, 'h21f8f, 'h21f8d, 'h10760, 'h108f2, 'h10770, 'h10780, 'h108f3, 'h10790, 'h10af0, 'h107a0, 'h108f4, 'h107b0, 'h107c0, 'h108f5, 'h107d0, 'h107e0, 'h108f6, 'h103bc, 'h107f0, 'h10800, 'h108f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10810, 'h10820, 'h108f8, 'h10830, 'h10840, 'h108f9, 'h10af0, 'h10850, 'h10860, 'h108fa, 'h10870, 'h10880, 'h108fb, 'h10890, 'h103bc, 'h108a0, 'h108fc, 'h108b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c0, 'h108fd, 'h108d0, 'h106e0, 'h108fe, 'h10b00, 'h106f0, 'h10700, 'h108ff, 'h10710, 'h10720, 'h10900, 'h10730, 'h10740, 'h10901, 'h103bc, 'h10750, 'h10760, 'h10902, 'h21f8e, 'h21f8f, 'h21f8d, 'h10770, 'h10780, 'h10903, 'h10790, 'h10b00, 'h107a0, 'h10904, 'h107b0, 'h107c0, 'h10905, 'h107d0, 'h107e0, 'h10906, 'h107f0, 'h103bc, 'h10800, 'h10907, 'h10810, 'h21f8e, 'h21f8f, 'h21f8d, 'h10820, 'h10908, 'h10830, 'h10840, 'h10909, 'h10b00, 'h10850, 'h10860, 'h1090a, 'h10870, 'h10880, 'h1090b, 'h10890, 'h108a0, 'h1090c, 'h103bc, 'h108b0, 'h108c0, 'h1090d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d0, 'h106e0, 'h1090e, 'h10b10, 'h106f0, 'h10700, 'h1090f, 'h10710, 'h10720, 'h10910, 'h10730, 'h10740, 'h10911, 'h10750, 'h103bc, 'h10760, 'h10912, 'h10770, 'h21f8e, 'h21f8f, 'h21f8d, 'h10780, 'h10913, 'h10790, 'h10b10, 'h107a0, 'h10914, 'h107b0, 'h107c0, 'h10915, 'h107d0, 'h107e0, 'h10916, 'h107f0, 'h10800, 'h10917, 'h103bc, 'h10810, 'h10820, 'h10918, 'h21f8e, 'h21f8f, 'h21f8d, 'h10830, 'h10840, 'h10919, 'h10b10, 'h10850, 'h10860, 'h1091a, 'h10870, 'h10880, 'h1091b, 'h10890, 'h108a0, 'h1091c, 'h108b0, 'h103bc, 'h108c0, 'h1091d, 'h108d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1091e, 'h10b20, 'h106f0, 'h10700, 'h1091f, 'h10710, 'h10720, 'h10920, 'h10730, 'h10740, 'h10921, 'h10750, 'h10760, 'h10922, 'h103bc, 'h10770, 'h10780, 'h10923, 'h21f8e, 'h21f8f, 'h21f8d, 'h10790, 'h10b20, 'h107a0, 'h10924, 'h107b0, 'h107c0, 'h10925, 'h107d0, 'h107e0, 'h10926, 'h107f0, 'h10800, 'h10927, 'h10810, 'h103bc, 'h10820, 'h10928, 'h10830, 'h21f8e, 'h21f8f, 'h21f8d, 'h10840, 'h10929, 'h10b20, 'h10850, 'h10860, 'h1092a, 'h10870, 'h10880, 'h1092b, 'h10890, 'h108a0, 'h1092c, 'h108b0, 'h108c0, 'h1092d, 'h103bc, 'h108d0, 'h106e0, 'h1092e, 'h10b30, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f0, 'h10700, 'h1092f, 'h10710, 'h10720, 'h10930, 'h10730, 'h10740, 'h10931, 'h10750, 'h10760, 'h10932, 'h10770, 'h103bc, 'h10780, 'h10933, 'h10790, 'h10b30, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a0, 'h10934, 'h107b0, 'h107c0, 'h10935, 'h107d0, 'h107e0, 'h10936, 'h107f0, 'h10800, 'h10937, 'h10810, 'h10820, 'h10938, 'h103bc, 'h10830, 'h10840, 'h10939, 'h10b30, 'h21f8e, 'h21f8f, 'h21f8d, 'h10850, 'h10860, 'h1093a, 'h10870, 'h10880, 'h1093b, 'h10890, 'h108a0, 'h1093c, 'h108b0, 'h108c0, 'h1093d, 'h108d0, 'h103bc, 'h106e0, 'h1093e, 'h10b40, 'h106f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10700, 'h1093f, 'h10710, 'h10720, 'h10940, 'h10730, 'h10740, 'h10941, 'h10750, 'h10760, 'h10942, 'h10770, 'h10780, 'h10943, 'h103bc, 'h10790, 'h10b40, 'h107a0, 'h10944, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b0, 'h107c0, 'h10945, 'h107d0, 'h107e0, 'h10946, 'h107f0, 'h10800, 'h10947, 'h10810, 'h10820, 'h10948, 'h10830, 'h103bc, 'h10840, 'h10949, 'h10b40, 'h10850, 'h21f8e, 'h21f8f, 'h21f8d, 'h10860, 'h1094a, 'h10870, 'h10880, 'h1094b, 'h10890, 'h108a0, 'h1094c, 'h108b0, 'h108c0, 'h1094d, 'h108d0, 'h106e0, 'h1094e, 'h10b50, 'h103bc, 'h106f0, 'h10700, 'h1094f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10710, 'h10720, 'h10950, 'h10730, 'h10740, 'h10951, 'h10750, 'h10760, 'h10952, 'h10770, 'h10780, 'h10953, 'h10790, 'h10b50, 'h103bc, 'h107a0, 'h10954, 'h107b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c0, 'h10955, 'h107d0, 'h107e0, 'h10956, 'h107f0, 'h10800, 'h10957, 'h10810, 'h10820, 'h10958, 'h10830, 'h10840, 'h10959, 'h10b50, 'h103bc, 'h10850, 'h10860, 'h1095a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10870, 'h10880, 'h1095b, 'h10890, 'h108a0, 'h1095c, 'h108b0, 'h108c0, 'h1095d, 'h108d0, 'h106e0, 'h1095e, 'h10b60, 'h106f0, 'h103bc, 'h10700, 'h1095f, 'h10710, 'h21f8e, 'h21f8f, 'h21f8d, 'h10720, 'h10960, 'h10730, 'h10740, 'h10961, 'h10750, 'h10760, 'h10962, 'h10770, 'h10780, 'h10963, 'h10790, 'h10b60, 'h107a0, 'h10964, 'h103bc, 'h107b0, 'h107c0, 'h10965, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d0, 'h107e0, 'h10966, 'h107f0, 'h10800, 'h10967, 'h10810, 'h10820, 'h10968, 'h10830, 'h10840, 'h10969, 'h10b60, 'h10850, 'h103bc, 'h10860, 'h1096a, 'h10870, 'h21f8e, 'h21f8f, 'h21f8d, 'h10880, 'h1096b, 'h10890, 'h108a0, 'h1096c, 'h108b0, 'h108c0, 'h1096d, 'h108d0, 'h106e0, 'h1096e, 'h10b70, 'h106f0, 'h10700, 'h1096f, 'h103bc, 'h10710, 'h10720, 'h10970, 'h21f8e, 'h21f8f, 'h21f8d, 'h10730, 'h10740, 'h10971, 'h10750, 'h10760, 'h10972, 'h10770, 'h10780, 'h10973, 'h10790, 'h10b70, 'h107a0, 'h10974, 'h107b0, 'h103bc, 'h107c0, 'h10975, 'h107d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e0, 'h10976, 'h107f0, 'h10800, 'h10977, 'h10810, 'h10820, 'h10978, 'h10830, 'h10840, 'h10979, 'h10b70, 'h10850, 'h10860, 'h1097a, 'h103bc, 'h10870, 'h10880, 'h1097b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10890, 'h108a0, 'h1097c, 'h108b0, 'h108c0, 'h1097d, 'h108d0, 'h106e0, 'h1097e, 'h10b80, 'h106f0, 'h10700, 'h1097f, 'h10710, 'h103bc, 'h10720, 'h10980, 'h10730, 'h21f8e, 'h21f8f, 'h21f8d, 'h10740, 'h10981, 'h10750, 'h10760, 'h10982, 'h10770, 'h10780, 'h10983, 'h10790, 'h10b80, 'h107a0, 'h10984, 'h107b0, 'h107c0, 'h10985, 'h103bc, 'h107d0, 'h107e0, 'h10986, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f0, 'h10800, 'h10987, 'h10810, 'h10820, 'h10988, 'h10830, 'h10840, 'h10989, 'h10b80, 'h10850, 'h10860, 'h1098a, 'h10870, 'h103bc, 'h10880, 'h1098b, 'h10890, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a0, 'h1098c, 'h108b0, 'h108c0, 'h1098d, 'h108d0, 'h106e0, 'h1098e, 'h10b90, 'h106f0, 'h10700, 'h1098f, 'h10710, 'h10720, 'h10990, 'h103bc, 'h10730, 'h10740, 'h10991, 'h21f8e, 'h21f8f, 'h21f8d, 'h10750, 'h10760, 'h10992, 'h10770, 'h10780, 'h10993, 'h10790, 'h10b90, 'h107a0, 'h10994, 'h107b0, 'h107c0, 'h10995, 'h107d0, 'h103bc, 'h107e0, 'h10996, 'h107f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10800, 'h10997, 'h10810, 'h10820, 'h10998, 'h10830, 'h10840, 'h10999, 'h10b90, 'h10850, 'h10860, 'h1099a, 'h10870, 'h10880, 'h1099b, 'h103bc, 'h10890, 'h108a0, 'h1099c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b0, 'h108c0, 'h1099d, 'h108d0, 'h106e0, 'h1099e, 'h10ba0, 'h106f0, 'h10700, 'h1099f, 'h10710, 'h10720, 'h109a0, 'h10730, 'h103bc, 'h10740, 'h109a1, 'h10750, 'h21f8e, 'h21f8f, 'h21f8d, 'h10760, 'h109a2, 'h10770, 'h10780, 'h109a3, 'h10790, 'h10ba0, 'h107a0, 'h109a4, 'h107b0, 'h107c0, 'h109a5, 'h107d0, 'h107e0, 'h109a6, 'h103bc, 'h107f0, 'h10800, 'h109a7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10810, 'h10820, 'h109a8, 'h10830, 'h10840, 'h109a9, 'h10ba0, 'h10850, 'h10860, 'h109aa, 'h10870, 'h10880, 'h109ab, 'h10890, 'h103bc, 'h108a0, 'h109ac, 'h108b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c0, 'h109ad, 'h108d0, 'h106e0, 'h109ae, 'h10bb0, 'h106f0, 'h10700, 'h109af, 'h10710, 'h10720, 'h109b0, 'h10730, 'h10740, 'h109b1, 'h103bc, 'h10750, 'h10760, 'h109b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10770, 'h10780, 'h109b3, 'h10790, 'h10bb0, 'h107a0, 'h109b4, 'h107b0, 'h107c0, 'h109b5, 'h107d0, 'h107e0, 'h109b6, 'h107f0, 'h103bc, 'h10800, 'h109b7, 'h10810, 'h21f8e, 'h21f8f, 'h21f8d, 'h10820, 'h109b8, 'h10830, 'h10840, 'h109b9, 'h10bb0, 'h10850, 'h10860, 'h109ba, 'h10870, 'h10880, 'h109bb, 'h10890, 'h108a0, 'h109bc, 'h103bc, 'h108b0, 'h108c0, 'h109bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d0, 'h106e0, 'h109be, 'h10bc0, 'h106f0, 'h10700, 'h109bf, 'h10710, 'h10720, 'h109c0, 'h10730, 'h10740, 'h109c1, 'h10750, 'h103bc, 'h10760, 'h109c2, 'h10770, 'h21f8e, 'h21f8f, 'h21f8d, 'h10780, 'h109c3, 'h10790, 'h10bc0, 'h107a0, 'h109c4, 'h107b0, 'h107c0, 'h109c5, 'h107d0, 'h107e0, 'h109c6, 'h107f0, 'h10800, 'h109c7, 'h103bc, 'h10810, 'h10820, 'h109c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10830, 'h10840, 'h109c9, 'h10bc0, 'h10850, 'h10860, 'h109ca, 'h10870, 'h10880, 'h109cb, 'h10890, 'h108a0, 'h109cc, 'h108b0, 'h103bc, 'h108c0, 'h109cd, 'h108d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h109ce, 'h10bd0, 'h106f0, 'h10700, 'h109cf, 'h10710, 'h10720, 'h109d0, 'h10730, 'h10740, 'h109d1, 'h10750, 'h10760, 'h109d2, 'h103bc, 'h10770, 'h10780, 'h109d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10790, 'h10bd0, 'h107a0, 'h109d4, 'h107b0, 'h107c0, 'h109d5, 'h107d0, 'h107e0, 'h109d6, 'h107f0, 'h10800, 'h109d7, 'h10810, 'h103bc, 'h10820, 'h109d8, 'h10830, 'h21f8e, 'h21f8f, 'h21f8d, 'h10840, 'h109d9, 'h10bd0, 'h10850, 'h10860, 'h109da, 'h10870, 'h10880, 'h109db, 'h10890, 'h108a0, 'h109dc, 'h108b0, 'h108c0, 'h109dd, 'h103bc, 'h108d0, 'h106e0, 'h109de, 'h10be0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f0, 'h10700, 'h109df, 'h10710, 'h10720, 'h109e0, 'h10730, 'h10740, 'h109e1, 'h10750, 'h10760, 'h109e2, 'h10770, 'h103bc, 'h10780, 'h109e3, 'h10790, 'h10be0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a0, 'h109e4, 'h107b0, 'h107c0, 'h109e5, 'h107d0, 'h107e0, 'h109e6, 'h107f0, 'h10800, 'h109e7, 'h10810, 'h10820, 'h109e8, 'h103bc, 'h10830, 'h10840, 'h109e9, 'h10be0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10850, 'h10860, 'h109ea, 'h10870, 'h10880, 'h109eb, 'h10890, 'h108a0, 'h109ec, 'h108b0, 'h108c0, 'h109ed, 'h108d0, 'h103bc, 'h106e0, 'h109ee, 'h10bf0, 'h106f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10700, 'h109ef, 'h10710, 'h10720, 'h109f0, 'h10730, 'h10740, 'h109f1, 'h10750, 'h10760, 'h109f2, 'h10770, 'h10780, 'h109f3, 'h103bc, 'h10790, 'h10bf0, 'h107a0, 'h109f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b0, 'h107c0, 'h109f5, 'h107d0, 'h107e0, 'h109f6, 'h107f0, 'h10800, 'h109f7, 'h10810, 'h10820, 'h109f8, 'h10830, 'h103bc, 'h10840, 'h109f9, 'h10bf0, 'h10850, 'h21f8e, 'h21f8f, 'h21f8d, 'h10860, 'h109fa, 'h10870, 'h10880, 'h109fb, 'h10890, 'h108a0, 'h109fc, 'h108b0, 'h108c0, 'h109fd, 'h108d0, 'h106e0, 'h109fe, 'h10c00, 'h103bc, 'h106f0, 'h10700, 'h109ff, 'h21f8e, 'h21f8f, 'h21f8d, 'h10710, 'h10720, 'h10a00, 'h10730, 'h10740, 'h10a01, 'h10750, 'h10760, 'h10a02, 'h10770, 'h10780, 'h10a03, 'h10790, 'h10c00, 'h103bc, 'h107a0, 'h10a04, 'h107b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c0, 'h10a05, 'h107d0, 'h107e0, 'h10a06, 'h107f0, 'h10800, 'h10a07, 'h10810, 'h10820, 'h10a08, 'h10830, 'h10840, 'h10a09, 'h10c00, 'h103bc, 'h10850, 'h10860, 'h10a0a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10870, 'h10880, 'h10a0b, 'h10890, 'h108a0, 'h10a0c, 'h108b0, 'h108c0, 'h10a0d, 'h108d0, 'h106e0, 'h10a0e, 'h10c10, 'h106f0, 'h103bc, 'h10700, 'h10a0f, 'h10710, 'h21f8e, 'h21f8f, 'h21f8d, 'h10720, 'h10a10, 'h10730, 'h10740, 'h10a11, 'h10750, 'h10760, 'h10a12, 'h10770, 'h10780, 'h10a13, 'h10790, 'h10c10, 'h107a0, 'h10a14, 'h103bc, 'h107b0, 'h107c0, 'h10a15, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d0, 'h107e0, 'h10a16, 'h107f0, 'h10800, 'h10a17, 'h10810, 'h10820, 'h10a18, 'h10830, 'h10840, 'h10a19, 'h10c10, 'h10850, 'h103bc, 'h10860, 'h10a1a, 'h10870, 'h21f8e, 'h21f8f, 'h21f8d, 'h10880, 'h10a1b, 'h10890, 'h108a0, 'h10a1c, 'h108b0, 'h108c0, 'h10a1d, 'h108d0, 'h106e0, 'h10a1e, 'h10c20, 'h106f0, 'h10700, 'h10a1f, 'h103bc, 'h10710, 'h10720, 'h10a20, 'h21f8e, 'h21f8f, 'h21f8d, 'h10730, 'h10740, 'h10a21, 'h10750, 'h10760, 'h10a22, 'h10770, 'h10780, 'h10a23, 'h10790, 'h10c20, 'h107a0, 'h10a24, 'h107b0, 'h103bc, 'h107c0, 'h10a25, 'h107d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e0, 'h10a26, 'h107f0, 'h10800, 'h10a27, 'h10810, 'h10820, 'h10a28, 'h10830, 'h10840, 'h10a29, 'h10c20, 'h10850, 'h10860, 'h10a2a, 'h103bc, 'h10870, 'h10880, 'h10a2b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10890, 'h108a0, 'h10a2c, 'h108b0, 'h108c0, 'h10a2d, 'h108d0, 'h106e0, 'h10a2e, 'h10c30, 'h106f0, 'h10700, 'h10a2f, 'h10710, 'h103bc, 'h10720, 'h10a30, 'h10730, 'h21f8e, 'h21f8f, 'h21f8d, 'h10740, 'h10a31, 'h10750, 'h10760, 'h10a32, 'h10770, 'h10780, 'h10a33, 'h10790, 'h10c30, 'h107a0, 'h10a34, 'h107b0, 'h107c0, 'h10a35, 'h103bc, 'h107d0, 'h107e0, 'h10a36, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f0, 'h10800, 'h10a37, 'h10810, 'h10820, 'h10a38, 'h10830, 'h10840, 'h10a39, 'h10c30, 'h10850, 'h10860, 'h10a3a, 'h10870, 'h103bc, 'h10880, 'h10a3b, 'h10890, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a0, 'h10a3c, 'h108b0, 'h108c0, 'h10a3d, 'h108d0, 'h106e0, 'h10a3e, 'h10c40, 'h106f0, 'h10700, 'h10a3f, 'h10710, 'h10720, 'h10a40, 'h103bc, 'h10730, 'h10740, 'h10a41, 'h21f8e, 'h21f8f, 'h21f8d, 'h10750, 'h10760, 'h10a42, 'h10770, 'h10780, 'h10a43, 'h10790, 'h10c40, 'h107a0, 'h10a44, 'h107b0, 'h107c0, 'h10a45, 'h107d0, 'h103bc, 'h107e0, 'h10a46, 'h107f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10800, 'h10a47, 'h10810, 'h10820, 'h10a48, 'h10830, 'h10840, 'h10a49, 'h10c40, 'h10850, 'h10860, 'h10a4a, 'h10870, 'h10880, 'h10a4b, 'h103bc, 'h10890, 'h108a0, 'h10a4c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b0, 'h108c0, 'h10a4d, 'h108d0, 'h106e0, 'h10a4e, 'h10c50, 'h106f0, 'h10700, 'h10a4f, 'h10710, 'h10720, 'h10a50, 'h10730, 'h103bc, 'h10740, 'h10a51, 'h10750, 'h21f8e, 'h21f8f, 'h21f8d, 'h10760, 'h10a52, 'h10770, 'h10780, 'h10a53, 'h10790, 'h10c50, 'h107a0, 'h10a54, 'h107b0, 'h107c0, 'h10a55, 'h107d0, 'h107e0, 'h10a56, 'h103bc, 'h107f0, 'h10800, 'h10a57, 'h21f8e, 'h21f8f, 'h21f8d, 'h10810, 'h10820, 'h10a58, 'h10830, 'h10840, 'h10a59, 'h10c50, 'h10850, 'h10860, 'h10a5a, 'h10870, 'h10880, 'h10a5b, 'h10890, 'h103bc, 'h108a0, 'h10a5c, 'h108b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c0, 'h10a5d, 'h108d0, 'h106e0, 'h10a5e, 'h10c60, 'h106f0, 'h10700, 'h10a5f, 'h10710, 'h10720, 'h10a60, 'h10730, 'h10740, 'h10a61, 'h103bc, 'h10750, 'h10760, 'h10a62, 'h21f8e, 'h21f8f, 'h21f8d, 'h10770, 'h10780, 'h10a63, 'h10790, 'h10c60, 'h107a0, 'h10a64, 'h107b0, 'h107c0, 'h10a65, 'h107d0, 'h107e0, 'h10a66, 'h107f0, 'h103bc, 'h10800, 'h10a67, 'h10810, 'h21f8e, 'h21f8f, 'h21f8d, 'h10820, 'h10a68, 'h10830, 'h10840, 'h10a69, 'h10c60, 'h10850, 'h10860, 'h10a6a, 'h10870, 'h10880, 'h10a6b, 'h10890, 'h108a0, 'h10a6c, 'h103bc, 'h108b0, 'h108c0, 'h10a6d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d0, 'h106e0, 'h10a6e, 'h10c70, 'h106f0, 'h10700, 'h10a6f, 'h10710, 'h10720, 'h10a70, 'h10730, 'h10740, 'h10a71, 'h10750, 'h103bc, 'h10760, 'h10a72, 'h10770, 'h21f8e, 'h21f8f, 'h21f8d, 'h10780, 'h10a73, 'h10790, 'h10c70, 'h107a0, 'h10a74, 'h107b0, 'h107c0, 'h10a75, 'h107d0, 'h107e0, 'h10a76, 'h107f0, 'h10800, 'h10a77, 'h103bc, 'h10810, 'h10820, 'h10a78, 'h21f8e, 'h21f8f, 'h21f8d, 'h10830, 'h10840, 'h10a79, 'h10c70, 'h10850, 'h10860, 'h10a7a, 'h10870, 'h10880, 'h10a7b, 'h10890, 'h108a0, 'h10a7c, 'h108b0, 'h103bc, 'h108c0, 'h10a7d, 'h108d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h10a7e, 'h10c80, 'h106f0, 'h10700, 'h10a7f, 'h10710, 'h10720, 'h10a80, 'h10730, 'h10740, 'h10a81, 'h10750, 'h10760, 'h10a82, 'h103bc, 'h10770, 'h10780, 'h10a83, 'h21f8e, 'h21f8f, 'h21f8d, 'h10790, 'h10c80, 'h107a0, 'h10a84, 'h107b0, 'h107c0, 'h10a85, 'h107d0, 'h107e0, 'h10a86, 'h107f0, 'h10800, 'h10a87, 'h10810, 'h103bc, 'h10820, 'h10a88, 'h10830, 'h21f8e, 'h21f8f, 'h21f8d, 'h10840, 'h10a89, 'h10c80, 'h10850, 'h10860, 'h10a8a, 'h10870, 'h10880, 'h10a8b, 'h10890, 'h108a0, 'h10a8c, 'h108b0, 'h108c0, 'h10a8d, 'h103bc, 'h108d0, 'h106e0, 'h10a8e, 'h10c90, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f0, 'h10700, 'h10a8f, 'h10710, 'h10720, 'h10a90, 'h10730, 'h10740, 'h10a91, 'h10750, 'h10760, 'h10a92, 'h10770, 'h103bc, 'h10780, 'h10a93, 'h10790, 'h10c90, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a0, 'h10a94, 'h107b0, 'h107c0, 'h10a95, 'h107d0, 'h107e0, 'h10a96, 'h107f0, 'h10800, 'h10a97, 'h10810, 'h10820, 'h10a98, 'h103bc, 'h10830, 'h10840, 'h10a99, 'h10c90, 'h21f8e, 'h21f8f, 'h21f8d, 'h10850, 'h10860, 'h10a9a, 'h10870, 'h10880, 'h10a9b, 'h10890, 'h108a0, 'h10a9c, 'h108b0, 'h108c0, 'h10a9d, 'h108d0, 'h103bc, 'h106e0, 'h10a9e, 'h10ca0, 'h106f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10700, 'h10a9f, 'h10710, 'h10720, 'h10aa0, 'h10730, 'h10740, 'h10aa1, 'h10750, 'h10760, 'h10aa2, 'h10770, 'h10780, 'h10aa3, 'h103bc, 'h10790, 'h10ca0, 'h107a0, 'h10aa4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b0, 'h107c0, 'h10aa5, 'h107d0, 'h107e0, 'h10aa6, 'h107f0, 'h10800, 'h10aa7, 'h10810, 'h10820, 'h10aa8, 'h10830, 'h103bc, 'h10840, 'h10aa9, 'h10ca0, 'h10850, 'h21f8e, 'h21f8f, 'h21f8d, 'h10860, 'h10aaa, 'h10870, 'h10880, 'h10aab, 'h10890, 'h108a0, 'h10aac, 'h108b0, 'h108c0, 'h10aad, 'h108d0, 'h106e0, 'h10aae, 'h10cb0, 'h103bc, 'h106f0, 'h10700, 'h10aaf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10710, 'h10720, 'h10ab0, 'h10730, 'h10740, 'h10ab1, 'h10750, 'h10760, 'h10ab2, 'h10770, 'h10780, 'h10ab3, 'h10790, 'h10cb0, 'h103bc, 'h107a0, 'h10ab4, 'h107b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c0, 'h10ab5, 'h107d0, 'h107e0, 'h10ab6, 'h107f0, 'h10800, 'h10ab7, 'h10810, 'h10820, 'h10ab8, 'h10830, 'h10840, 'h10ab9, 'h10cb0, 'h103bc, 'h10850, 'h10860, 'h10aba, 'h21f8e, 'h21f8f, 'h21f8d, 'h10870, 'h10880, 'h10abb, 'h10890, 'h108a0, 'h10abc, 'h108b0, 'h108c0, 'h10abd, 'h108d0, 'h106e0, 'h10abe, 'h10cc0, 'h106f0, 'h103bc, 'h10700, 'h10abf, 'h10710, 'h21f8e, 'h21f8f, 'h21f8d, 'h10720, 'h10ac0, 'h10730, 'h10740, 'h10ac1, 'h10750, 'h10760, 'h10ac2, 'h10770, 'h10780, 'h10ac3, 'h10790, 'h10cc0, 'h107a0, 'h10ac4, 'h103bc, 'h107b0, 'h107c0, 'h10ac5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d0, 'h107e0, 'h10ac6, 'h107f0, 'h10800, 'h10ac7, 'h10810, 'h10820, 'h10ac8, 'h10830, 'h10840, 'h10ac9, 'h10cc0, 'h10850, 'h103bc, 'h10860, 'h10aca, 'h10870, 'h21f8e, 'h21f8f, 'h21f8d, 'h10880, 'h10acb, 'h10890, 'h108a0, 'h10acc, 'h108b0, 'h108c0, 'h10acd, 'h108d0, 'h106e0, 'h10ace, 'h10cd0, 'h106f0, 'h10700, 'h10acf, 'h103bc, 'h10710, 'h10720, 'h10ad0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10730, 'h10740, 'h10ad1, 'h10750, 'h10760, 'h10ad2, 'h10770, 'h10780, 'h10ad3, 'h10790, 'h10cd0, 'h107a0, 'h10ad4, 'h107b0, 'h103bc, 'h107c0, 'h10ad5, 'h107d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e0, 'h10ad6, 'h107f0, 'h10800, 'h10ad7, 'h10810, 'h10820, 'h10ad8, 'h10830, 'h10840, 'h10ad9, 'h10cd0, 'h10850, 'h10860, 'h10ada, 'h103bc, 'h10870, 'h10880, 'h10adb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10890, 'h108a0, 'h10adc, 'h108b0, 'h108c0, 'h10add, 'h108d0, 'h106e0, 'h108de, 'h10ae0, 'h106f0, 'h10700, 'h108df, 'h10710, 'h103bc, 'h10720, 'h108e0, 'h10730, 'h21f8e, 'h21f8f, 'h21f8d, 'h10740, 'h108e1, 'h10750, 'h10760, 'h108e2, 'h10770, 'h10780, 'h108e3, 'h10790, 'h10ae0, 'h107a0, 'h108e4, 'h107b0, 'h107c0, 'h108e5, 'h103bc, 'h107d0, 'h107e0, 'h108e6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f0, 'h10800, 'h108e7, 'h10810, 'h10820, 'h108e8, 'h10830, 'h10840, 'h108e9, 'h10ae0, 'h10850, 'h10860, 'h108ea, 'h10870, 'h103bc, 'h10880, 'h108eb, 'h10890, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a0, 'h108ec, 'h108b0, 'h108c0, 'h108ed, 'h108d0, 'h106e0, 'h108ee, 'h10af0, 'h106f0, 'h10700, 'h108ef, 'h10710, 'h10720, 'h108f0, 'h103bc, 'h10730, 'h10740, 'h108f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10750, 'h10760, 'h108f2, 'h10770, 'h10780, 'h108f3, 'h10790, 'h10af0, 'h107a0, 'h108f4, 'h107b0, 'h107c0, 'h108f5, 'h107d0, 'h103bc, 'h107e0, 'h108f6, 'h107f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10800, 'h108f7, 'h10810, 'h10820, 'h108f8, 'h10830, 'h10840, 'h108f9, 'h10af0, 'h10850, 'h10860, 'h108fa, 'h10870, 'h10880, 'h108fb, 'h103bc, 'h10890, 'h108a0, 'h108fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b0, 'h108c0, 'h108fd, 'h108d0, 'h106e0, 'h108fe, 'h10b00, 'h106f0, 'h10700, 'h108ff, 'h10710, 'h10720, 'h10900, 'h10730, 'h103bc, 'h10740, 'h10901, 'h10750, 'h21f8e, 'h21f8f, 'h21f8d, 'h10760, 'h10902, 'h10770, 'h10780, 'h10903, 'h10790, 'h10b00, 'h107a0, 'h10904, 'h107b0, 'h107c0, 'h10905, 'h107d0, 'h107e0, 'h10906, 'h103bc, 'h107f0, 'h10800, 'h10907, 'h21f8e, 'h21f8f, 'h21f8d, 'h10810, 'h10820, 'h10908, 'h10830, 'h10840, 'h10909, 'h10b00, 'h10850, 'h10860, 'h1090a, 'h10870, 'h10880, 'h1090b, 'h10890, 'h103bc, 'h108a0, 'h1090c, 'h108b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c0, 'h1090d, 'h108d0, 'h106e0, 'h1090e, 'h10b10, 'h106f0, 'h10700, 'h1090f, 'h10710, 'h10720, 'h10910, 'h10730, 'h10740, 'h10911, 'h103bc, 'h10750, 'h10760, 'h10912, 'h21f8e, 'h21f8f, 'h21f8d, 'h10770, 'h10780, 'h10913, 'h10790, 'h10b10, 'h107a0, 'h10914, 'h107b0, 'h107c0, 'h10915, 'h107d0, 'h107e0, 'h10916, 'h107f0, 'h103bc, 'h10800, 'h10917, 'h10810, 'h21f8e, 'h21f8f, 'h21f8d, 'h10820, 'h10918, 'h10830, 'h10840, 'h10919, 'h10b10, 'h10850, 'h10860, 'h1091a, 'h10870, 'h10880, 'h1091b, 'h10890, 'h108a0, 'h1091c, 'h103bc, 'h108b0, 'h108c0, 'h1091d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d0, 'h106e0, 'h1091e, 'h10b20, 'h106f0, 'h10700, 'h1091f, 'h10710, 'h10720, 'h10920, 'h10730, 'h10740, 'h10921, 'h10750, 'h103bc, 'h10760, 'h10922, 'h10770, 'h21f8e, 'h21f8f, 'h21f8d, 'h10780, 'h10923, 'h10790, 'h10b20, 'h107a0, 'h10924, 'h107b0, 'h107c0, 'h10925, 'h107d0, 'h107e0, 'h10926, 'h107f0, 'h10800, 'h10927, 'h103bc, 'h10810, 'h10820, 'h10928, 'h21f8e, 'h21f8f, 'h21f8d, 'h10830, 'h10840, 'h10929, 'h10b20, 'h10850, 'h10860, 'h1092a, 'h10870, 'h10880, 'h1092b, 'h10890, 'h108a0, 'h1092c, 'h108b0, 'h103bc, 'h108c0, 'h1092d, 'h108d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1092e, 'h10b30, 'h106f0, 'h10700, 'h1092f, 'h10710, 'h10720, 'h10930, 'h10730, 'h10740, 'h10931, 'h10750, 'h10760, 'h10932, 'h103bc, 'h10770, 'h10780, 'h10933, 'h21f8e, 'h21f8f, 'h21f8d, 'h10790, 'h10b30, 'h107a0, 'h10934, 'h107b0, 'h107c0, 'h10935, 'h107d0, 'h107e0, 'h10936, 'h107f0, 'h10800, 'h10937, 'h10810, 'h103bc, 'h10820, 'h10938, 'h10830, 'h21f8e, 'h21f8f, 'h21f8d, 'h10840, 'h10939, 'h10b30, 'h10850, 'h10860, 'h1093a, 'h10870, 'h10880, 'h1093b, 'h10890, 'h108a0, 'h1093c, 'h108b0, 'h108c0, 'h1093d, 'h103bc, 'h108d0, 'h106e0, 'h1093e, 'h10b40, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f0, 'h10700, 'h1093f, 'h10710, 'h10720, 'h10940, 'h10730, 'h10740, 'h10941, 'h10750, 'h10760, 'h10942, 'h10770, 'h103bc, 'h10780, 'h10943, 'h10790, 'h10b40, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a0, 'h10944, 'h107b0, 'h107c0, 'h10945, 'h107d0, 'h107e0, 'h10946, 'h107f0, 'h10800, 'h10947, 'h10810, 'h10820, 'h10948, 'h103bc, 'h10830, 'h10840, 'h10949, 'h10b40, 'h21f8e, 'h21f8f, 'h21f8d, 'h10850, 'h10860, 'h1094a, 'h10870, 'h10880, 'h1094b, 'h10890, 'h108a0, 'h1094c, 'h108b0, 'h108c0, 'h1094d, 'h108d0, 'h103bc, 'h106e0, 'h1094e, 'h10b50, 'h106f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10700, 'h1094f, 'h10710, 'h10720, 'h10950, 'h10730, 'h10740, 'h10951, 'h10750, 'h10760, 'h10952, 'h10770, 'h10780, 'h10953, 'h103bc, 'h10790, 'h10b50, 'h107a0, 'h10954, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b0, 'h107c0, 'h10955, 'h107d0, 'h107e0, 'h10956, 'h107f0, 'h10800, 'h10957, 'h10810, 'h10820, 'h10958, 'h10830, 'h103bc, 'h10840, 'h10959, 'h10b50, 'h10850, 'h21f8e, 'h21f8f, 'h21f8d, 'h10860, 'h1095a, 'h10870, 'h10880, 'h1095b, 'h10890, 'h108a0, 'h1095c, 'h108b0, 'h108c0, 'h1095d, 'h108d0, 'h106e0, 'h1095e, 'h10b60, 'h103bc, 'h106f0, 'h10700, 'h1095f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10710, 'h10720, 'h10960, 'h10730, 'h10740, 'h10961, 'h10750, 'h10760, 'h10962, 'h10770, 'h10780, 'h10963, 'h10790, 'h10b60, 'h103bc, 'h107a0, 'h10964, 'h107b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c0, 'h10965, 'h107d0, 'h107e0, 'h10966, 'h107f0, 'h10800, 'h10967, 'h10810, 'h10820, 'h10968, 'h10830, 'h10840, 'h10969, 'h10b60, 'h103bc, 'h10850, 'h10860, 'h1096a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10870, 'h10880, 'h1096b, 'h10890, 'h108a0, 'h1096c, 'h108b0, 'h108c0, 'h1096d, 'h108d0, 'h106e0, 'h1096e, 'h10b70, 'h106f0, 'h103bc, 'h10700, 'h1096f, 'h10710, 'h21f8e, 'h21f8f, 'h21f8d, 'h10720, 'h10970, 'h10730, 'h10740, 'h10971, 'h10750, 'h10760, 'h10972, 'h10770, 'h10780, 'h10973, 'h10790, 'h10b70, 'h107a0, 'h10974, 'h103bc, 'h107b0, 'h107c0, 'h10975, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d0, 'h107e0, 'h10976, 'h107f0, 'h10800, 'h10977, 'h10810, 'h10820, 'h10978, 'h10830, 'h10840, 'h10979, 'h10b70, 'h10850, 'h103bc, 'h10860, 'h1097a, 'h10870, 'h21f8e, 'h21f8f, 'h21f8d, 'h10880, 'h1097b, 'h10890, 'h108a0, 'h1097c, 'h108b0, 'h108c0, 'h1097d, 'h108d0, 'h106e0, 'h1097e, 'h10b80, 'h106f0, 'h10700, 'h1097f, 'h103bc, 'h10710, 'h10720, 'h10980, 'h21f8e, 'h21f8f, 'h21f8d, 'h10730, 'h10740, 'h10981, 'h10750, 'h10760, 'h10982, 'h10770, 'h10780, 'h10983, 'h10790, 'h10b80, 'h107a0, 'h10984, 'h107b0, 'h103bc, 'h107c0, 'h10985, 'h107d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e0, 'h10986, 'h107f0, 'h10800, 'h10987, 'h10810, 'h10820, 'h10988, 'h10830, 'h10840, 'h10989, 'h10b80, 'h10850, 'h10860, 'h1098a, 'h103bc, 'h10870, 'h10880, 'h1098b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10890, 'h108a0, 'h1098c, 'h108b0, 'h108c0, 'h1098d, 'h108d0, 'h106e0, 'h1098e, 'h10b90, 'h106f0, 'h10700, 'h1098f, 'h10710, 'h103bc, 'h10720, 'h10990, 'h10730, 'h21f8e, 'h21f8f, 'h21f8d, 'h10740, 'h10991, 'h10750, 'h10760, 'h10992, 'h10770, 'h10780, 'h10993, 'h10790, 'h10b90, 'h107a0, 'h10994, 'h107b0, 'h107c0, 'h10995, 'h103bc, 'h107d0, 'h107e0, 'h10996, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f0, 'h10800, 'h10997, 'h10810, 'h10820, 'h10998, 'h10830, 'h10840, 'h10999, 'h10b90, 'h10850, 'h10860, 'h1099a, 'h10870, 'h103bc, 'h10880, 'h1099b, 'h10890, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a0, 'h1099c, 'h108b0, 'h108c0, 'h1099d, 'h108d0, 'h106e0, 'h1099e, 'h10ba0, 'h106f0, 'h10700, 'h1099f, 'h10710, 'h10720, 'h109a0, 'h103bc, 'h10730, 'h10740, 'h109a1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10750, 'h10760, 'h109a2, 'h10770, 'h10780, 'h109a3, 'h10790, 'h10ba0, 'h107a0, 'h109a4, 'h107b0, 'h107c0, 'h109a5, 'h107d0, 'h103bc, 'h107e0, 'h109a6, 'h107f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10800, 'h109a7, 'h10810, 'h10820, 'h109a8, 'h10830, 'h10840, 'h109a9, 'h10ba0, 'h10850, 'h10860, 'h109aa, 'h10870, 'h10880, 'h109ab, 'h103bc, 'h10890, 'h108a0, 'h109ac, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b0, 'h108c0, 'h109ad, 'h108d0, 'h106e0, 'h109ae, 'h10bb0, 'h106f0, 'h10700, 'h109af, 'h10710, 'h10720, 'h109b0, 'h10730, 'h103bc, 'h10740, 'h109b1, 'h10750, 'h21f8e, 'h21f8f, 'h21f8d, 'h10760, 'h109b2, 'h10770, 'h10780, 'h109b3, 'h10790, 'h10bb0, 'h107a0, 'h109b4, 'h107b0, 'h107c0, 'h109b5, 'h107d0, 'h107e0, 'h109b6, 'h103bc, 'h107f0, 'h10800, 'h109b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10810, 'h10820, 'h109b8, 'h10830, 'h10840, 'h109b9, 'h10bb0, 'h10850, 'h10860, 'h109ba, 'h10870, 'h10880, 'h109bb, 'h10890, 'h103bc, 'h108a0, 'h109bc, 'h108b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c0, 'h109bd, 'h108d0, 'h106e0, 'h109be, 'h10bc0, 'h106f0, 'h10700, 'h109bf, 'h10710, 'h10720, 'h109c0, 'h10730, 'h10740, 'h109c1, 'h103bc, 'h10750, 'h10760, 'h109c2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10770, 'h10780, 'h109c3, 'h10790, 'h10bc0, 'h107a0, 'h109c4, 'h107b0, 'h107c0, 'h109c5, 'h107d0, 'h107e0, 'h109c6, 'h107f0, 'h103bc, 'h10800, 'h109c7, 'h10810, 'h21f8e, 'h21f8f, 'h21f8d, 'h10820, 'h109c8, 'h10830, 'h10840, 'h109c9, 'h10bc0, 'h10850, 'h10860, 'h109ca, 'h10870, 'h10880, 'h109cb, 'h10890, 'h108a0, 'h109cc, 'h103bc, 'h108b0, 'h108c0, 'h109cd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d0, 'h106e0, 'h109ce, 'h10bd0, 'h106f0, 'h10700, 'h109cf, 'h10710, 'h10720, 'h109d0, 'h10730, 'h10740, 'h109d1, 'h10750, 'h103bc, 'h10760, 'h109d2, 'h10770, 'h21f8e, 'h21f8f, 'h21f8d, 'h10780, 'h109d3, 'h10790, 'h10bd0, 'h107a0, 'h109d4, 'h107b0, 'h107c0, 'h109d5, 'h107d0, 'h107e0, 'h109d6, 'h107f0, 'h10800, 'h109d7, 'h103bc, 'h10810, 'h10820, 'h109d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10830, 'h10840, 'h109d9, 'h10bd0, 'h10850, 'h10860, 'h109da, 'h10870, 'h10880, 'h109db, 'h10890, 'h108a0, 'h109dc, 'h108b0, 'h103bc, 'h108c0, 'h109dd, 'h108d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h109de, 'h10be0, 'h106f0, 'h10700, 'h109df, 'h10710, 'h10720, 'h109e0, 'h10730, 'h10740, 'h109e1, 'h10750, 'h10760, 'h109e2, 'h103bc, 'h10770, 'h10780, 'h109e3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10790, 'h10be0, 'h107a0, 'h109e4, 'h107b0, 'h107c0, 'h109e5, 'h107d0, 'h107e0, 'h109e6, 'h107f0, 'h10800, 'h109e7, 'h10810, 'h103bc, 'h10820, 'h109e8, 'h10830, 'h21f8e, 'h21f8f, 'h21f8d, 'h10840, 'h109e9, 'h10be0, 'h10850, 'h10860, 'h109ea, 'h10870, 'h10880, 'h109eb, 'h10890, 'h108a0, 'h109ec, 'h108b0, 'h108c0, 'h109ed, 'h103bc, 'h108d0, 'h106e0, 'h109ee, 'h10bf0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f0, 'h10700, 'h109ef, 'h10710, 'h10720, 'h109f0, 'h10730, 'h10740, 'h109f1, 'h10750, 'h10760, 'h109f2, 'h10770, 'h103bc, 'h10780, 'h109f3, 'h10790, 'h10bf0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a0, 'h109f4, 'h107b0, 'h107c0, 'h109f5, 'h107d0, 'h107e0, 'h109f6, 'h107f0, 'h10800, 'h109f7, 'h10810, 'h10820, 'h109f8, 'h103bc, 'h10830, 'h10840, 'h109f9, 'h10bf0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10850, 'h10860, 'h109fa, 'h10870, 'h10880, 'h109fb, 'h10890, 'h108a0, 'h109fc, 'h108b0, 'h108c0, 'h109fd, 'h108d0, 'h103bc, 'h106e0, 'h109fe, 'h10c00, 'h106f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10700, 'h109ff, 'h10710, 'h10720, 'h10a00, 'h10730, 'h10740, 'h10a01, 'h10750, 'h10760, 'h10a02, 'h10770, 'h10780, 'h10a03, 'h103bc, 'h10790, 'h10c00, 'h107a0, 'h10a04, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b0, 'h107c0, 'h10a05, 'h107d0, 'h107e0, 'h10a06, 'h107f0, 'h10800, 'h10a07, 'h10810, 'h10820, 'h10a08, 'h10830, 'h103bc, 'h10840, 'h10a09, 'h10c00, 'h10850, 'h21f8e, 'h21f8f, 'h21f8d, 'h10860, 'h10a0a, 'h10870, 'h10880, 'h10a0b, 'h10890, 'h108a0, 'h10a0c, 'h108b0, 'h108c0, 'h10a0d, 'h108d0, 'h106e0, 'h10a0e, 'h10c10, 'h103bc, 'h106f0, 'h10700, 'h10a0f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10710, 'h10720, 'h10a10, 'h10730, 'h10740, 'h10a11, 'h10750, 'h10760, 'h10a12, 'h10770, 'h10780, 'h10a13, 'h10790, 'h10c10, 'h103bc, 'h107a0, 'h10a14, 'h107b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c0, 'h10a15, 'h107d0, 'h107e0, 'h10a16, 'h107f0, 'h10800, 'h10a17, 'h10810, 'h10820, 'h10a18, 'h10830, 'h10840, 'h10a19, 'h10c10, 'h103bc, 'h10850, 'h10860, 'h10a1a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10870, 'h10880, 'h10a1b, 'h10890, 'h108a0, 'h10a1c, 'h108b0, 'h108c0, 'h10a1d, 'h108d0, 'h106e0, 'h10a1e, 'h10c20, 'h106f0, 'h103bc, 'h10700, 'h10a1f, 'h10710, 'h21f8e, 'h21f8f, 'h21f8d, 'h10720, 'h10a20, 'h10730, 'h10740, 'h10a21, 'h10750, 'h10760, 'h10a22, 'h10770, 'h10780, 'h10a23, 'h10790, 'h10c20, 'h107a0, 'h10a24, 'h103bc, 'h107b0, 'h107c0, 'h10a25, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d0, 'h107e0, 'h10a26, 'h107f0, 'h10800, 'h10a27, 'h10810, 'h10820, 'h10a28, 'h10830, 'h10840, 'h10a29, 'h10c20, 'h10850, 'h103bc, 'h10860, 'h10a2a, 'h10870, 'h21f8e, 'h21f8f, 'h21f8d, 'h10880, 'h10a2b, 'h10890, 'h108a0, 'h10a2c, 'h108b0, 'h108c0, 'h10a2d, 'h108d0, 'h106e0, 'h10a2e, 'h10c30, 'h106f0, 'h10700, 'h10a2f, 'h103bc, 'h10710, 'h10720, 'h10a30, 'h21f8e, 'h21f8f, 'h21f8d, 'h10730, 'h10740, 'h10a31, 'h10750, 'h10760, 'h10a32, 'h10770, 'h10780, 'h10a33, 'h10790, 'h10c30, 'h107a0, 'h10a34, 'h107b0, 'h103bc, 'h107c0, 'h10a35, 'h107d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e0, 'h10a36, 'h107f0, 'h10800, 'h10a37, 'h10810, 'h10820, 'h10a38, 'h10830, 'h10840, 'h10a39, 'h10c30, 'h10850, 'h10860, 'h10a3a, 'h103bc, 'h10870, 'h10880, 'h10a3b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10890, 'h108a0, 'h10a3c, 'h108b0, 'h108c0, 'h10a3d, 'h108d0, 'h106e0, 'h10a3e, 'h10c40, 'h106f0, 'h10700, 'h10a3f, 'h10710, 'h103bc, 'h10720, 'h10a40, 'h10730, 'h21f8e, 'h21f8f, 'h21f8d, 'h10740, 'h10a41, 'h10750, 'h10760, 'h10a42, 'h10770, 'h10780, 'h10a43, 'h10790, 'h10c40, 'h107a0, 'h10a44, 'h107b0, 'h107c0, 'h10a45, 'h103bc, 'h107d0, 'h107e0, 'h10a46, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f0, 'h10800, 'h10a47, 'h10810, 'h10820, 'h10a48, 'h10830, 'h10840, 'h10a49, 'h10c40, 'h10850, 'h10860, 'h10a4a, 'h10870, 'h103bc, 'h10880, 'h10a4b, 'h10890, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a0, 'h10a4c, 'h108b0, 'h108c0, 'h10a4d, 'h108d0, 'h106e0, 'h10a4e, 'h10c50, 'h106f0, 'h10700, 'h10a4f, 'h10710, 'h10720, 'h10a50, 'h103bc, 'h10730, 'h10740, 'h10a51, 'h21f8e, 'h21f8f, 'h21f8d, 'h10750, 'h10760, 'h10a52, 'h10770, 'h10780, 'h10a53, 'h10790, 'h10c50, 'h107a0, 'h10a54, 'h107b0, 'h107c0, 'h10a55, 'h107d0, 'h103bc, 'h107e0, 'h10a56, 'h107f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10800, 'h10a57, 'h10810, 'h10820, 'h10a58, 'h10830, 'h10840, 'h10a59, 'h10c50, 'h10850, 'h10860, 'h10a5a, 'h10870, 'h10880, 'h10a5b, 'h103bc, 'h10890, 'h108a0, 'h10a5c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b0, 'h108c0, 'h10a5d, 'h108d0, 'h106e0, 'h10a5e, 'h10c60, 'h106f0, 'h10700, 'h10a5f, 'h10710, 'h10720, 'h10a60, 'h10730, 'h103bc, 'h10740, 'h10a61, 'h10750, 'h21f8e, 'h21f8f, 'h21f8d, 'h10760, 'h10a62, 'h10770, 'h10780, 'h10a63, 'h10790, 'h10c60, 'h107a0, 'h10a64, 'h107b0, 'h107c0, 'h10a65, 'h107d0, 'h107e0, 'h10a66, 'h103bc, 'h107f0, 'h10800, 'h10a67, 'h21f8e, 'h21f8f, 'h21f8d, 'h10810, 'h10820, 'h10a68, 'h10830, 'h10840, 'h10a69, 'h10c60, 'h10850, 'h10860, 'h10a6a, 'h10870, 'h10880, 'h10a6b, 'h10890, 'h103bc, 'h108a0, 'h10a6c, 'h108b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c0, 'h10a6d, 'h108d0, 'h106e0, 'h10a6e, 'h10c70, 'h106f0, 'h10700, 'h10a6f, 'h10710, 'h10720, 'h10a70, 'h10730, 'h10740, 'h10a71, 'h103bc, 'h10750, 'h10760, 'h10a72, 'h21f8e, 'h21f8f, 'h21f8d, 'h10770, 'h10780, 'h10a73, 'h10790, 'h10c70, 'h107a0, 'h10a74, 'h107b0, 'h107c0, 'h10a75, 'h107d0, 'h107e0, 'h10a76, 'h107f0, 'h103bc, 'h10800, 'h10a77, 'h10810, 'h21f8e, 'h21f8f, 'h21f8d, 'h10820, 'h10a78, 'h10830, 'h10840, 'h10a79, 'h10c70, 'h10850, 'h10860, 'h10a7a, 'h10870, 'h10880, 'h10a7b, 'h10890, 'h108a0, 'h10a7c, 'h103bc, 'h108b0, 'h108c0, 'h10a7d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d0, 'h106e0, 'h10a7e, 'h10c80, 'h106f0, 'h10700, 'h10a7f, 'h10710, 'h10720, 'h10a80, 'h10730, 'h10740, 'h10a81, 'h10750, 'h103bc, 'h10760, 'h10a82, 'h10770, 'h21f8e, 'h21f8f, 'h21f8d, 'h10780, 'h10a83, 'h10790, 'h10c80, 'h107a0, 'h10a84, 'h107b0, 'h107c0, 'h10a85, 'h107d0, 'h107e0, 'h10a86, 'h107f0, 'h10800, 'h10a87, 'h103bc, 'h10810, 'h10820, 'h10a88, 'h21f8e, 'h21f8f, 'h21f8d, 'h10830, 'h10840, 'h10a89, 'h10c80, 'h10850, 'h10860, 'h10a8a, 'h10870, 'h10880, 'h10a8b, 'h10890, 'h108a0, 'h10a8c, 'h108b0, 'h103bc, 'h108c0, 'h10a8d, 'h108d0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h10a8e, 'h10c90, 'h106f0, 'h10700, 'h10a8f, 'h10710, 'h10720, 'h10a90, 'h10730, 'h10740, 'h10a91, 'h10750, 'h10760, 'h10a92, 'h103bc, 'h10770, 'h10780, 'h10a93, 'h21f8e, 'h21f8f, 'h21f8d, 'h10790, 'h10c90, 'h107a0, 'h10a94, 'h107b0, 'h107c0, 'h10a95, 'h107d0, 'h107e0, 'h10a96, 'h107f0, 'h10800, 'h10a97, 'h10810, 'h103bc, 'h10820, 'h10a98, 'h10830, 'h21f8e, 'h21f8f, 'h21f8d, 'h10840, 'h10a99, 'h10c90, 'h10850, 'h10860, 'h10a9a, 'h10870, 'h10880, 'h10a9b, 'h10890, 'h108a0, 'h10a9c, 'h108b0, 'h108c0, 'h10a9d, 'h103bc, 'h108d0, 'h106e0, 'h10a9e, 'h10ca0, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f0, 'h10700, 'h10a9f, 'h10710, 'h10720, 'h10aa0, 'h10730, 'h10740, 'h10aa1, 'h10750, 'h10760, 'h10aa2, 'h10770, 'h103bc, 'h10780, 'h10aa3, 'h10790, 'h10ca0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a0, 'h10aa4, 'h107b0, 'h107c0, 'h10aa5, 'h107d0, 'h107e0, 'h10aa6, 'h107f0, 'h10800, 'h10aa7, 'h10810, 'h10820, 'h10aa8, 'h103bc, 'h10830, 'h10840, 'h10aa9, 'h10ca0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10850, 'h10860, 'h10aaa, 'h10870, 'h10880, 'h10aab, 'h10890, 'h108a0, 'h10aac, 'h108b0, 'h108c0, 'h10aad, 'h108d0, 'h103bc, 'h106e0, 'h10aae, 'h10cb0, 'h106f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10700, 'h10aaf, 'h10710, 'h10720, 'h10ab0, 'h10730, 'h10740, 'h10ab1, 'h10750, 'h10760, 'h10ab2, 'h10770, 'h10780, 'h10ab3, 'h103bc, 'h10790, 'h10cb0, 'h107a0, 'h10ab4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b0, 'h107c0, 'h10ab5, 'h107d0, 'h107e0, 'h10ab6, 'h107f0, 'h10800, 'h10ab7, 'h10810, 'h10820, 'h10ab8, 'h10830, 'h103bc, 'h10840, 'h10ab9, 'h10cb0, 'h10850, 'h21f8e, 'h21f8f, 'h21f8d, 'h10860, 'h10aba, 'h10870, 'h10880, 'h10abb, 'h10890, 'h108a0, 'h10abc, 'h108b0, 'h108c0, 'h10abd, 'h108d0, 'h106e0, 'h10abe, 'h10cc0, 'h103bc, 'h106f0, 'h10700, 'h10abf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10710, 'h10720, 'h10ac0, 'h10730, 'h10740, 'h10ac1, 'h10750, 'h10760, 'h10ac2, 'h10770, 'h10780, 'h10ac3, 'h10790, 'h10cc0, 'h103bc, 'h107a0, 'h10ac4, 'h107b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c0, 'h10ac5, 'h107d0, 'h107e0, 'h10ac6, 'h107f0, 'h10800, 'h10ac7, 'h10810, 'h10820, 'h10ac8, 'h10830, 'h10840, 'h10ac9, 'h10cc0, 'h103bc, 'h10850, 'h10860, 'h10aca, 'h21f8e, 'h21f8f, 'h21f8d, 'h10870, 'h10880, 'h10acb, 'h10890, 'h108a0, 'h10acc, 'h108b0, 'h108c0, 'h10acd, 'h108d0, 'h106e0, 'h10ace, 'h10cd0, 'h106f0, 'h103bc, 'h10700, 'h10acf, 'h10710, 'h21f8e, 'h21f8f, 'h21f8d, 'h10720, 'h10ad0, 'h10730, 'h10740, 'h10ad1, 'h10750, 'h10760, 'h10ad2, 'h10770, 'h10780, 'h10ad3, 'h10790, 'h10cd0, 'h107a0, 'h10ad4, 'h103bc, 'h107b0, 'h107c0, 'h10ad5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d0, 'h107e0, 'h10ad6, 'h107f0, 'h10800, 'h10ad7, 'h10810, 'h10820, 'h10ad8, 'h10830, 'h10840, 'h10ad9, 'h10cd0, 'h10850, 'h103bc, 'h10860, 'h10ada, 'h10870, 'h21f8e, 'h21f8f, 'h21f8d, 'h10880, 'h10adb, 'h10890, 'h108a0, 'h10adc, 'h108b0, 'h108c0, 'h10add, 'h108d0, 'h106e1, 'h108de, 'h10ae1, 'h106f1, 'h10701, 'h108df, 'h103bc, 'h10711, 'h10721, 'h108e0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10731, 'h10741, 'h108e1, 'h10751, 'h10761, 'h108e2, 'h10771, 'h10781, 'h108e3, 'h10791, 'h10ae1, 'h107a1, 'h108e4, 'h107b1, 'h103bc, 'h107c1, 'h108e5, 'h107d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e1, 'h108e6, 'h107f1, 'h10801, 'h108e7, 'h10811, 'h10821, 'h108e8, 'h10831, 'h10841, 'h108e9, 'h10ae1, 'h10851, 'h10861, 'h108ea, 'h103bc, 'h10871, 'h10881, 'h108eb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10891, 'h108a1, 'h108ec, 'h108b1, 'h108c1, 'h108ed, 'h108d1, 'h106e1, 'h108ee, 'h10af1, 'h106f1, 'h10701, 'h108ef, 'h10711, 'h103bc, 'h10721, 'h108f0, 'h10731, 'h21f8e, 'h21f8f, 'h21f8d, 'h10741, 'h108f1, 'h10751, 'h10761, 'h108f2, 'h10771, 'h10781, 'h108f3, 'h10791, 'h10af1, 'h107a1, 'h108f4, 'h107b1, 'h107c1, 'h108f5, 'h103bc, 'h107d1, 'h107e1, 'h108f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f1, 'h10801, 'h108f7, 'h10811, 'h10821, 'h108f8, 'h10831, 'h10841, 'h108f9, 'h10af1, 'h10851, 'h10861, 'h108fa, 'h10871, 'h103bc, 'h10881, 'h108fb, 'h10891, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a1, 'h108fc, 'h108b1, 'h108c1, 'h108fd, 'h108d1, 'h106e1, 'h108fe, 'h10b01, 'h106f1, 'h10701, 'h108ff, 'h10711, 'h10721, 'h10900, 'h103bc, 'h10731, 'h10741, 'h10901, 'h21f8e, 'h21f8f, 'h21f8d, 'h10751, 'h10761, 'h10902, 'h10771, 'h10781, 'h10903, 'h10791, 'h10b01, 'h107a1, 'h10904, 'h107b1, 'h107c1, 'h10905, 'h107d1, 'h103bc, 'h107e1, 'h10906, 'h107f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10801, 'h10907, 'h10811, 'h10821, 'h10908, 'h10831, 'h10841, 'h10909, 'h10b01, 'h10851, 'h10861, 'h1090a, 'h10871, 'h10881, 'h1090b, 'h103bc, 'h10891, 'h108a1, 'h1090c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b1, 'h108c1, 'h1090d, 'h108d1, 'h106e1, 'h1090e, 'h10b11, 'h106f1, 'h10701, 'h1090f, 'h10711, 'h10721, 'h10910, 'h10731, 'h103bc, 'h10741, 'h10911, 'h10751, 'h21f8e, 'h21f8f, 'h21f8d, 'h10761, 'h10912, 'h10771, 'h10781, 'h10913, 'h10791, 'h10b11, 'h107a1, 'h10914, 'h107b1, 'h107c1, 'h10915, 'h107d1, 'h107e1, 'h10916, 'h103bc, 'h107f1, 'h10801, 'h10917, 'h21f8e, 'h21f8f, 'h21f8d, 'h10811, 'h10821, 'h10918, 'h10831, 'h10841, 'h10919, 'h10b11, 'h10851, 'h10861, 'h1091a, 'h10871, 'h10881, 'h1091b, 'h10891, 'h103bc, 'h108a1, 'h1091c, 'h108b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c1, 'h1091d, 'h108d1, 'h106e1, 'h1091e, 'h10b21, 'h106f1, 'h10701, 'h1091f, 'h10711, 'h10721, 'h10920, 'h10731, 'h10741, 'h10921, 'h103bc, 'h10751, 'h10761, 'h10922, 'h21f8e, 'h21f8f, 'h21f8d, 'h10771, 'h10781, 'h10923, 'h10791, 'h10b21, 'h107a1, 'h10924, 'h107b1, 'h107c1, 'h10925, 'h107d1, 'h107e1, 'h10926, 'h107f1, 'h103bc, 'h10801, 'h10927, 'h10811, 'h21f8e, 'h21f8f, 'h21f8d, 'h10821, 'h10928, 'h10831, 'h10841, 'h10929, 'h10b21, 'h10851, 'h10861, 'h1092a, 'h10871, 'h10881, 'h1092b, 'h10891, 'h108a1, 'h1092c, 'h103bc, 'h108b1, 'h108c1, 'h1092d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d1, 'h106e1, 'h1092e, 'h10b31, 'h106f1, 'h10701, 'h1092f, 'h10711, 'h10721, 'h10930, 'h10731, 'h10741, 'h10931, 'h10751, 'h103bc, 'h10761, 'h10932, 'h10771, 'h21f8e, 'h21f8f, 'h21f8d, 'h10781, 'h10933, 'h10791, 'h10b31, 'h107a1, 'h10934, 'h107b1, 'h107c1, 'h10935, 'h107d1, 'h107e1, 'h10936, 'h107f1, 'h10801, 'h10937, 'h103bc, 'h10811, 'h10821, 'h10938, 'h21f8e, 'h21f8f, 'h21f8d, 'h10831, 'h10841, 'h10939, 'h10b31, 'h10851, 'h10861, 'h1093a, 'h10871, 'h10881, 'h1093b, 'h10891, 'h108a1, 'h1093c, 'h108b1, 'h103bc, 'h108c1, 'h1093d, 'h108d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1093e, 'h10b41, 'h106f1, 'h10701, 'h1093f, 'h10711, 'h10721, 'h10940, 'h10731, 'h10741, 'h10941, 'h10751, 'h10761, 'h10942, 'h103bc, 'h10771, 'h10781, 'h10943, 'h21f8e, 'h21f8f, 'h21f8d, 'h10791, 'h10b41, 'h107a1, 'h10944, 'h107b1, 'h107c1, 'h10945, 'h107d1, 'h107e1, 'h10946, 'h107f1, 'h10801, 'h10947, 'h10811, 'h103bc, 'h10821, 'h10948, 'h10831, 'h21f8e, 'h21f8f, 'h21f8d, 'h10841, 'h10949, 'h10b41, 'h10851, 'h10861, 'h1094a, 'h10871, 'h10881, 'h1094b, 'h10891, 'h108a1, 'h1094c, 'h108b1, 'h108c1, 'h1094d, 'h103bc, 'h108d1, 'h106e1, 'h1094e, 'h10b51, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f1, 'h10701, 'h1094f, 'h10711, 'h10721, 'h10950, 'h10731, 'h10741, 'h10951, 'h10751, 'h10761, 'h10952, 'h10771, 'h103bc, 'h10781, 'h10953, 'h10791, 'h10b51, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a1, 'h10954, 'h107b1, 'h107c1, 'h10955, 'h107d1, 'h107e1, 'h10956, 'h107f1, 'h10801, 'h10957, 'h10811, 'h10821, 'h10958, 'h103bc, 'h10831, 'h10841, 'h10959, 'h10b51, 'h21f8e, 'h21f8f, 'h21f8d, 'h10851, 'h10861, 'h1095a, 'h10871, 'h10881, 'h1095b, 'h10891, 'h108a1, 'h1095c, 'h108b1, 'h108c1, 'h1095d, 'h108d1, 'h103bc, 'h106e1, 'h1095e, 'h10b61, 'h106f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10701, 'h1095f, 'h10711, 'h10721, 'h10960, 'h10731, 'h10741, 'h10961, 'h10751, 'h10761, 'h10962, 'h10771, 'h10781, 'h10963, 'h103bc, 'h10791, 'h10b61, 'h107a1, 'h10964, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b1, 'h107c1, 'h10965, 'h107d1, 'h107e1, 'h10966, 'h107f1, 'h10801, 'h10967, 'h10811, 'h10821, 'h10968, 'h10831, 'h103bc, 'h10841, 'h10969, 'h10b61, 'h10851, 'h21f8e, 'h21f8f, 'h21f8d, 'h10861, 'h1096a, 'h10871, 'h10881, 'h1096b, 'h10891, 'h108a1, 'h1096c, 'h108b1, 'h108c1, 'h1096d, 'h108d1, 'h106e1, 'h1096e, 'h10b71, 'h103bc, 'h106f1, 'h10701, 'h1096f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10711, 'h10721, 'h10970, 'h10731, 'h10741, 'h10971, 'h10751, 'h10761, 'h10972, 'h10771, 'h10781, 'h10973, 'h10791, 'h10b71, 'h103bc, 'h107a1, 'h10974, 'h107b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c1, 'h10975, 'h107d1, 'h107e1, 'h10976, 'h107f1, 'h10801, 'h10977, 'h10811, 'h10821, 'h10978, 'h10831, 'h10841, 'h10979, 'h10b71, 'h103bc, 'h10851, 'h10861, 'h1097a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10871, 'h10881, 'h1097b, 'h10891, 'h108a1, 'h1097c, 'h108b1, 'h108c1, 'h1097d, 'h108d1, 'h106e1, 'h1097e, 'h10b81, 'h106f1, 'h103bc, 'h10701, 'h1097f, 'h10711, 'h21f8e, 'h21f8f, 'h21f8d, 'h10721, 'h10980, 'h10731, 'h10741, 'h10981, 'h10751, 'h10761, 'h10982, 'h10771, 'h10781, 'h10983, 'h10791, 'h10b81, 'h107a1, 'h10984, 'h103bc, 'h107b1, 'h107c1, 'h10985, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d1, 'h107e1, 'h10986, 'h107f1, 'h10801, 'h10987, 'h10811, 'h10821, 'h10988, 'h10831, 'h10841, 'h10989, 'h10b81, 'h10851, 'h103bc, 'h10861, 'h1098a, 'h10871, 'h21f8e, 'h21f8f, 'h21f8d, 'h10881, 'h1098b, 'h10891, 'h108a1, 'h1098c, 'h108b1, 'h108c1, 'h1098d, 'h108d1, 'h106e1, 'h1098e, 'h10b91, 'h106f1, 'h10701, 'h1098f, 'h103bc, 'h10711, 'h10721, 'h10990, 'h21f8e, 'h21f8f, 'h21f8d, 'h10731, 'h10741, 'h10991, 'h10751, 'h10761, 'h10992, 'h10771, 'h10781, 'h10993, 'h10791, 'h10b91, 'h107a1, 'h10994, 'h107b1, 'h103bc, 'h107c1, 'h10995, 'h107d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e1, 'h10996, 'h107f1, 'h10801, 'h10997, 'h10811, 'h10821, 'h10998, 'h10831, 'h10841, 'h10999, 'h10b91, 'h10851, 'h10861, 'h1099a, 'h103bc, 'h10871, 'h10881, 'h1099b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10891, 'h108a1, 'h1099c, 'h108b1, 'h108c1, 'h1099d, 'h108d1, 'h106e1, 'h1099e, 'h10ba1, 'h106f1, 'h10701, 'h1099f, 'h10711, 'h103bc, 'h10721, 'h109a0, 'h10731, 'h21f8e, 'h21f8f, 'h21f8d, 'h10741, 'h109a1, 'h10751, 'h10761, 'h109a2, 'h10771, 'h10781, 'h109a3, 'h10791, 'h10ba1, 'h107a1, 'h109a4, 'h107b1, 'h107c1, 'h109a5, 'h103bc, 'h107d1, 'h107e1, 'h109a6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f1, 'h10801, 'h109a7, 'h10811, 'h10821, 'h109a8, 'h10831, 'h10841, 'h109a9, 'h10ba1, 'h10851, 'h10861, 'h109aa, 'h10871, 'h103bc, 'h10881, 'h109ab, 'h10891, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a1, 'h109ac, 'h108b1, 'h108c1, 'h109ad, 'h108d1, 'h106e1, 'h109ae, 'h10bb1, 'h106f1, 'h10701, 'h109af, 'h10711, 'h10721, 'h109b0, 'h103bc, 'h10731, 'h10741, 'h109b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10751, 'h10761, 'h109b2, 'h10771, 'h10781, 'h109b3, 'h10791, 'h10bb1, 'h107a1, 'h109b4, 'h107b1, 'h107c1, 'h109b5, 'h107d1, 'h103bc, 'h107e1, 'h109b6, 'h107f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10801, 'h109b7, 'h10811, 'h10821, 'h109b8, 'h10831, 'h10841, 'h109b9, 'h10bb1, 'h10851, 'h10861, 'h109ba, 'h10871, 'h10881, 'h109bb, 'h103bc, 'h10891, 'h108a1, 'h109bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b1, 'h108c1, 'h109bd, 'h108d1, 'h106e1, 'h109be, 'h10bc1, 'h106f1, 'h10701, 'h109bf, 'h10711, 'h10721, 'h109c0, 'h10731, 'h103bc, 'h10741, 'h109c1, 'h10751, 'h21f8e, 'h21f8f, 'h21f8d, 'h10761, 'h109c2, 'h10771, 'h10781, 'h109c3, 'h10791, 'h10bc1, 'h107a1, 'h109c4, 'h107b1, 'h107c1, 'h109c5, 'h107d1, 'h107e1, 'h109c6, 'h103bc, 'h107f1, 'h10801, 'h109c7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10811, 'h10821, 'h109c8, 'h10831, 'h10841, 'h109c9, 'h10bc1, 'h10851, 'h10861, 'h109ca, 'h10871, 'h10881, 'h109cb, 'h10891, 'h103bc, 'h108a1, 'h109cc, 'h108b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c1, 'h109cd, 'h108d1, 'h106e1, 'h109ce, 'h10bd1, 'h106f1, 'h10701, 'h109cf, 'h10711, 'h10721, 'h109d0, 'h10731, 'h10741, 'h109d1, 'h103bc, 'h10751, 'h10761, 'h109d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10771, 'h10781, 'h109d3, 'h10791, 'h10bd1, 'h107a1, 'h109d4, 'h107b1, 'h107c1, 'h109d5, 'h107d1, 'h107e1, 'h109d6, 'h107f1, 'h103bc, 'h10801, 'h109d7, 'h10811, 'h21f8e, 'h21f8f, 'h21f8d, 'h10821, 'h109d8, 'h10831, 'h10841, 'h109d9, 'h10bd1, 'h10851, 'h10861, 'h109da, 'h10871, 'h10881, 'h109db, 'h10891, 'h108a1, 'h109dc, 'h103bc, 'h108b1, 'h108c1, 'h109dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d1, 'h106e1, 'h109de, 'h10be1, 'h106f1, 'h10701, 'h109df, 'h10711, 'h10721, 'h109e0, 'h10731, 'h10741, 'h109e1, 'h10751, 'h103bc, 'h10761, 'h109e2, 'h10771, 'h21f8e, 'h21f8f, 'h21f8d, 'h10781, 'h109e3, 'h10791, 'h10be1, 'h107a1, 'h109e4, 'h107b1, 'h107c1, 'h109e5, 'h107d1, 'h107e1, 'h109e6, 'h107f1, 'h10801, 'h109e7, 'h103bc, 'h10811, 'h10821, 'h109e8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10831, 'h10841, 'h109e9, 'h10be1, 'h10851, 'h10861, 'h109ea, 'h10871, 'h10881, 'h109eb, 'h10891, 'h108a1, 'h109ec, 'h108b1, 'h103bc, 'h108c1, 'h109ed, 'h108d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h109ee, 'h10bf1, 'h106f1, 'h10701, 'h109ef, 'h10711, 'h10721, 'h109f0, 'h10731, 'h10741, 'h109f1, 'h10751, 'h10761, 'h109f2, 'h103bc, 'h10771, 'h10781, 'h109f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10791, 'h10bf1, 'h107a1, 'h109f4, 'h107b1, 'h107c1, 'h109f5, 'h107d1, 'h107e1, 'h109f6, 'h107f1, 'h10801, 'h109f7, 'h10811, 'h103bc, 'h10821, 'h109f8, 'h10831, 'h21f8e, 'h21f8f, 'h21f8d, 'h10841, 'h109f9, 'h10bf1, 'h10851, 'h10861, 'h109fa, 'h10871, 'h10881, 'h109fb, 'h10891, 'h108a1, 'h109fc, 'h108b1, 'h108c1, 'h109fd, 'h103bc, 'h108d1, 'h106e1, 'h109fe, 'h10c01, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f1, 'h10701, 'h109ff, 'h10711, 'h10721, 'h10a00, 'h10731, 'h10741, 'h10a01, 'h10751, 'h10761, 'h10a02, 'h10771, 'h103bc, 'h10781, 'h10a03, 'h10791, 'h10c01, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a1, 'h10a04, 'h107b1, 'h107c1, 'h10a05, 'h107d1, 'h107e1, 'h10a06, 'h107f1, 'h10801, 'h10a07, 'h10811, 'h10821, 'h10a08, 'h103bc, 'h10831, 'h10841, 'h10a09, 'h10c01, 'h21f8e, 'h21f8f, 'h21f8d, 'h10851, 'h10861, 'h10a0a, 'h10871, 'h10881, 'h10a0b, 'h10891, 'h108a1, 'h10a0c, 'h108b1, 'h108c1, 'h10a0d, 'h108d1, 'h103bc, 'h106e1, 'h10a0e, 'h10c11, 'h106f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10701, 'h10a0f, 'h10711, 'h10721, 'h10a10, 'h10731, 'h10741, 'h10a11, 'h10751, 'h10761, 'h10a12, 'h10771, 'h10781, 'h10a13, 'h103bc, 'h10791, 'h10c11, 'h107a1, 'h10a14, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b1, 'h107c1, 'h10a15, 'h107d1, 'h107e1, 'h10a16, 'h107f1, 'h10801, 'h10a17, 'h10811, 'h10821, 'h10a18, 'h10831, 'h103bc, 'h10841, 'h10a19, 'h10c11, 'h10851, 'h21f8e, 'h21f8f, 'h21f8d, 'h10861, 'h10a1a, 'h10871, 'h10881, 'h10a1b, 'h10891, 'h108a1, 'h10a1c, 'h108b1, 'h108c1, 'h10a1d, 'h108d1, 'h106e1, 'h10a1e, 'h10c21, 'h103bc, 'h106f1, 'h10701, 'h10a1f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10711, 'h10721, 'h10a20, 'h10731, 'h10741, 'h10a21, 'h10751, 'h10761, 'h10a22, 'h10771, 'h10781, 'h10a23, 'h10791, 'h10c21, 'h103bc, 'h107a1, 'h10a24, 'h107b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c1, 'h10a25, 'h107d1, 'h107e1, 'h10a26, 'h107f1, 'h10801, 'h10a27, 'h10811, 'h10821, 'h10a28, 'h10831, 'h10841, 'h10a29, 'h10c21, 'h103bc, 'h10851, 'h10861, 'h10a2a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10871, 'h10881, 'h10a2b, 'h10891, 'h108a1, 'h10a2c, 'h108b1, 'h108c1, 'h10a2d, 'h108d1, 'h106e1, 'h10a2e, 'h10c31, 'h106f1, 'h103bc, 'h10701, 'h10a2f, 'h10711, 'h21f8e, 'h21f8f, 'h21f8d, 'h10721, 'h10a30, 'h10731, 'h10741, 'h10a31, 'h10751, 'h10761, 'h10a32, 'h10771, 'h10781, 'h10a33, 'h10791, 'h10c31, 'h107a1, 'h10a34, 'h103bc, 'h107b1, 'h107c1, 'h10a35, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d1, 'h107e1, 'h10a36, 'h107f1, 'h10801, 'h10a37, 'h10811, 'h10821, 'h10a38, 'h10831, 'h10841, 'h10a39, 'h10c31, 'h10851, 'h103bc, 'h10861, 'h10a3a, 'h10871, 'h21f8e, 'h21f8f, 'h21f8d, 'h10881, 'h10a3b, 'h10891, 'h108a1, 'h10a3c, 'h108b1, 'h108c1, 'h10a3d, 'h108d1, 'h106e1, 'h10a3e, 'h10c41, 'h106f1, 'h10701, 'h10a3f, 'h103bc, 'h10711, 'h10721, 'h10a40, 'h21f8e, 'h21f8f, 'h21f8d, 'h10731, 'h10741, 'h10a41, 'h10751, 'h10761, 'h10a42, 'h10771, 'h10781, 'h10a43, 'h10791, 'h10c41, 'h107a1, 'h10a44, 'h107b1, 'h103bc, 'h107c1, 'h10a45, 'h107d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e1, 'h10a46, 'h107f1, 'h10801, 'h10a47, 'h10811, 'h10821, 'h10a48, 'h10831, 'h10841, 'h10a49, 'h10c41, 'h10851, 'h10861, 'h10a4a, 'h103bc, 'h10871, 'h10881, 'h10a4b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10891, 'h108a1, 'h10a4c, 'h108b1, 'h108c1, 'h10a4d, 'h108d1, 'h106e1, 'h10a4e, 'h10c51, 'h106f1, 'h10701, 'h10a4f, 'h10711, 'h103bc, 'h10721, 'h10a50, 'h10731, 'h21f8e, 'h21f8f, 'h21f8d, 'h10741, 'h10a51, 'h10751, 'h10761, 'h10a52, 'h10771, 'h10781, 'h10a53, 'h10791, 'h10c51, 'h107a1, 'h10a54, 'h107b1, 'h107c1, 'h10a55, 'h103bc, 'h107d1, 'h107e1, 'h10a56, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f1, 'h10801, 'h10a57, 'h10811, 'h10821, 'h10a58, 'h10831, 'h10841, 'h10a59, 'h10c51, 'h10851, 'h10861, 'h10a5a, 'h10871, 'h103bc, 'h10881, 'h10a5b, 'h10891, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a1, 'h10a5c, 'h108b1, 'h108c1, 'h10a5d, 'h108d1, 'h106e1, 'h10a5e, 'h10c61, 'h106f1, 'h10701, 'h10a5f, 'h10711, 'h10721, 'h10a60, 'h103bc, 'h10731, 'h10741, 'h10a61, 'h21f8e, 'h21f8f, 'h21f8d, 'h10751, 'h10761, 'h10a62, 'h10771, 'h10781, 'h10a63, 'h10791, 'h10c61, 'h107a1, 'h10a64, 'h107b1, 'h107c1, 'h10a65, 'h107d1, 'h103bc, 'h107e1, 'h10a66, 'h107f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10801, 'h10a67, 'h10811, 'h10821, 'h10a68, 'h10831, 'h10841, 'h10a69, 'h10c61, 'h10851, 'h10861, 'h10a6a, 'h10871, 'h10881, 'h10a6b, 'h103bc, 'h10891, 'h108a1, 'h10a6c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b1, 'h108c1, 'h10a6d, 'h108d1, 'h106e1, 'h10a6e, 'h10c71, 'h106f1, 'h10701, 'h10a6f, 'h10711, 'h10721, 'h10a70, 'h10731, 'h103bc, 'h10741, 'h10a71, 'h10751, 'h21f8e, 'h21f8f, 'h21f8d, 'h10761, 'h10a72, 'h10771, 'h10781, 'h10a73, 'h10791, 'h10c71, 'h107a1, 'h10a74, 'h107b1, 'h107c1, 'h10a75, 'h107d1, 'h107e1, 'h10a76, 'h103bc, 'h107f1, 'h10801, 'h10a77, 'h21f8e, 'h21f8f, 'h21f8d, 'h10811, 'h10821, 'h10a78, 'h10831, 'h10841, 'h10a79, 'h10c71, 'h10851, 'h10861, 'h10a7a, 'h10871, 'h10881, 'h10a7b, 'h10891, 'h103bc, 'h108a1, 'h10a7c, 'h108b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c1, 'h10a7d, 'h108d1, 'h106e1, 'h10a7e, 'h10c81, 'h106f1, 'h10701, 'h10a7f, 'h10711, 'h10721, 'h10a80, 'h10731, 'h10741, 'h10a81, 'h103bc, 'h10751, 'h10761, 'h10a82, 'h21f8e, 'h21f8f, 'h21f8d, 'h10771, 'h10781, 'h10a83, 'h10791, 'h10c81, 'h107a1, 'h10a84, 'h107b1, 'h107c1, 'h10a85, 'h107d1, 'h107e1, 'h10a86, 'h107f1, 'h103bc, 'h10801, 'h10a87, 'h10811, 'h21f8e, 'h21f8f, 'h21f8d, 'h10821, 'h10a88, 'h10831, 'h10841, 'h10a89, 'h10c81, 'h10851, 'h10861, 'h10a8a, 'h10871, 'h10881, 'h10a8b, 'h10891, 'h108a1, 'h10a8c, 'h103bc, 'h108b1, 'h108c1, 'h10a8d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d1, 'h106e1, 'h10a8e, 'h10c91, 'h106f1, 'h10701, 'h10a8f, 'h10711, 'h10721, 'h10a90, 'h10731, 'h10741, 'h10a91, 'h10751, 'h103bc, 'h10761, 'h10a92, 'h10771, 'h21f8e, 'h21f8f, 'h21f8d, 'h10781, 'h10a93, 'h10791, 'h10c91, 'h107a1, 'h10a94, 'h107b1, 'h107c1, 'h10a95, 'h107d1, 'h107e1, 'h10a96, 'h107f1, 'h10801, 'h10a97, 'h103bc, 'h10811, 'h10821, 'h10a98, 'h21f8e, 'h21f8f, 'h21f8d, 'h10831, 'h10841, 'h10a99, 'h10c91, 'h10851, 'h10861, 'h10a9a, 'h10871, 'h10881, 'h10a9b, 'h10891, 'h108a1, 'h10a9c, 'h108b1, 'h103bc, 'h108c1, 'h10a9d, 'h108d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h10a9e, 'h10ca1, 'h106f1, 'h10701, 'h10a9f, 'h10711, 'h10721, 'h10aa0, 'h10731, 'h10741, 'h10aa1, 'h10751, 'h10761, 'h10aa2, 'h103bc, 'h10771, 'h10781, 'h10aa3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10791, 'h10ca1, 'h107a1, 'h10aa4, 'h107b1, 'h107c1, 'h10aa5, 'h107d1, 'h107e1, 'h10aa6, 'h107f1, 'h10801, 'h10aa7, 'h10811, 'h103bc, 'h10821, 'h10aa8, 'h10831, 'h21f8e, 'h21f8f, 'h21f8d, 'h10841, 'h10aa9, 'h10ca1, 'h10851, 'h10861, 'h10aaa, 'h10871, 'h10881, 'h10aab, 'h10891, 'h108a1, 'h10aac, 'h108b1, 'h108c1, 'h10aad, 'h103bc, 'h108d1, 'h106e1, 'h10aae, 'h10cb1, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f1, 'h10701, 'h10aaf, 'h10711, 'h10721, 'h10ab0, 'h10731, 'h10741, 'h10ab1, 'h10751, 'h10761, 'h10ab2, 'h10771, 'h103bc, 'h10781, 'h10ab3, 'h10791, 'h10cb1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a1, 'h10ab4, 'h107b1, 'h107c1, 'h10ab5, 'h107d1, 'h107e1, 'h10ab6, 'h107f1, 'h10801, 'h10ab7, 'h10811, 'h10821, 'h10ab8, 'h103bc, 'h10831, 'h10841, 'h10ab9, 'h10cb1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10851, 'h10861, 'h10aba, 'h10871, 'h10881, 'h10abb, 'h10891, 'h108a1, 'h10abc, 'h108b1, 'h108c1, 'h10abd, 'h108d1, 'h103bc, 'h106e1, 'h10abe, 'h10cc1, 'h106f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10701, 'h10abf, 'h10711, 'h10721, 'h10ac0, 'h10731, 'h10741, 'h10ac1, 'h10751, 'h10761, 'h10ac2, 'h10771, 'h10781, 'h10ac3, 'h103bc, 'h10791, 'h10cc1, 'h107a1, 'h10ac4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b1, 'h107c1, 'h10ac5, 'h107d1, 'h107e1, 'h10ac6, 'h107f1, 'h10801, 'h10ac7, 'h10811, 'h10821, 'h10ac8, 'h10831, 'h103bc, 'h10841, 'h10ac9, 'h10cc1, 'h10851, 'h21f8e, 'h21f8f, 'h21f8d, 'h10861, 'h10aca, 'h10871, 'h10881, 'h10acb, 'h10891, 'h108a1, 'h10acc, 'h108b1, 'h108c1, 'h10acd, 'h108d1, 'h106e1, 'h10ace, 'h10cd1, 'h103bc, 'h106f1, 'h10701, 'h10acf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10711, 'h10721, 'h10ad0, 'h10731, 'h10741, 'h10ad1, 'h10751, 'h10761, 'h10ad2, 'h10771, 'h10781, 'h10ad3, 'h10791, 'h10cd1, 'h103bc, 'h107a1, 'h10ad4, 'h107b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c1, 'h10ad5, 'h107d1, 'h107e1, 'h10ad6, 'h107f1, 'h10801, 'h10ad7, 'h10811, 'h10821, 'h10ad8, 'h10831, 'h10841, 'h10ad9, 'h10cd1, 'h103bc, 'h10851, 'h10861, 'h10ada, 'h21f8e, 'h21f8f, 'h21f8d, 'h10871, 'h10881, 'h10adb};
	int DATA2 [2*SIZE-1:0] = {DATA1, DATA0};
	
endpackage
