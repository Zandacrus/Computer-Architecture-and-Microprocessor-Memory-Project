

package LU_PKG_1;
	
	parameter SIZE = 8500;
	
	int DATA1 [SIZE-1:0] = {'h2004f8, 'h10003c, 'h10006c, 'h2004f7, 'h1004f9, 'h100000, 'h100047, 'h100044, 'h10006e, 'h10006f, 'h100070, 'h100071, 'h100072, 'h100073, 'h100074, 'h100075, 'h100076, 'h100077, 'h100078, 'h100079, 'h10007a, 'h10007b, 'h10003c, 'h10007c, 'h2004f7, 'h10007d, 'h100000, 'h100047, 'h100044, 'h10007e, 'h10007f, 'h100080, 'h100081, 'h100082, 'h100083, 'h100084, 'h100085, 'h100086, 'h100087, 'h100088, 'h100089, 'h10008a, 'h10008b, 'h10003c, 'h10008c, 'h2004f7, 'h10008d, 'h100000, 'h100047, 'h100044, 'h10008e, 'h10008f, 'h100090, 'h100091, 'h100092, 'h100093, 'h100094, 'h100095, 'h100096, 'h100097, 'h100098, 'h100099, 'h10009a, 'h10009b, 'h10003c, 'h10009c, 'h2004f7, 'h10009d, 'h100000, 'h100047, 'h100044, 'h10009e, 'h10009f, 'h1000a0, 'h1000a1, 'h1000a2, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h1000a7, 'h1000a8, 'h1000a9, 'h1000aa, 'h1000ab, 'h10003c, 'h1000ac, 'h2004f7, 'h1000ad, 'h100000, 'h100047, 'h100044, 'h1000ae, 'h1000af, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h1000b7, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h10003c, 'h1000bc, 'h2004f7, 'h1000bd, 'h100000, 'h100047, 'h100044, 'h1000be, 'h1000bf, 'h1000c0, 'h1000c1, 'h1000c2, 'h1000c3, 'h1000c4, 'h1000c5, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h10003c, 'h1000cc, 'h2004f7, 'h1000cd, 'h100000, 'h100047, 'h100044, 'h1000ce, 'h1000cf, 'h1000d0, 'h1000d1, 'h1000d2, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h10003c, 'h1000dc, 'h2004f7, 'h1000dd, 'h100000, 'h100047, 'h100044, 'h1000de, 'h1000df, 'h1000e0, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h10003c, 'h1000ec, 'h2004f7, 'h1000ed, 'h100000, 'h100047, 'h100044, 'h1000ee, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h10003c, 'h1000fc, 'h2004f7, 'h1000fd, 'h100000, 'h100047, 'h100044, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10003c, 'h10010c, 'h2004f7, 'h10010d, 'h100000, 'h100047, 'h100044, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10003c, 'h10011c, 'h2004f7, 'h10011d, 'h100000, 'h100047, 'h100044, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10003c, 'h10012c, 'h2004f7, 'h10012d, 'h100000, 'h100047, 'h100044, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10003c, 'h10013c, 'h2004f7, 'h10013d, 'h100000, 'h100047, 'h100044, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10003c, 'h10014c, 'h2004f7, 'h10014d, 'h100000, 'h100047, 'h100044, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10003c, 'h10015c, 'h2004f7, 'h10015d, 'h100000, 'h100047, 'h100044, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10003c, 'h10016c, 'h2004f7, 'h10016d, 'h100000, 'h100047, 'h100044, 'h10016e, 'h10016f, 'h100170, 'h100171, 'h100172, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10003c, 'h10017c, 'h2004f7, 'h10017d, 'h100000, 'h100047, 'h100044, 'h10017e, 'h10017f, 'h100180, 'h100181, 'h100182, 'h100183, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10003c, 'h10018c, 'h2004f7, 'h10018d, 'h100000, 'h100047, 'h100044, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h100192, 'h100193, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h10019c, 'h2004f7, 'h10019d, 'h100000, 'h100047, 'h100044, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h10003c, 'h1001ac, 'h2004f7, 'h1001ad, 'h100000, 'h100047, 'h100044, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h10003c, 'h1001bc, 'h2004f7, 'h1001bd, 'h100000, 'h100047, 'h100044, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h10003c, 'h1001cc, 'h2004f7, 'h1001cd, 'h100000, 'h100047, 'h100044, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h10003c, 'h1001dc, 'h2004f7, 'h1001dd, 'h100000, 'h100047, 'h100044, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h10003c, 'h1001ec, 'h2004f7, 'h1001ed, 'h100000, 'h100047, 'h100044, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h10003c, 'h1001fc, 'h2004f7, 'h1001fd, 'h100000, 'h100047, 'h100044, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10003c, 'h10020c, 'h2004f7, 'h10020d, 'h100000, 'h100047, 'h100044, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100213, 'h100214, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10003c, 'h10021c, 'h2004f7, 'h10021d, 'h100000, 'h100047, 'h100044, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h100223, 'h100224, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10003c, 'h10022c, 'h2004f7, 'h10022d, 'h100000, 'h100047, 'h100044, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10003c, 'h10023c, 'h2004f7, 'h10023d, 'h100000, 'h100047, 'h100044, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10003c, 'h10024c, 'h2004f7, 'h10024d, 'h100000, 'h100047, 'h100044, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10003c, 'h10025c, 'h2004f7, 'h10025d, 'h100000, 'h100047, 'h100044, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10003c, 'h10026c, 'h2004f7, 'h10026d, 'h100000, 'h100047, 'h100044, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h2004f8, 'h10006e, 'h10006f, 'h100070, 'h100071, 'h100072, 'h100076, 'h100073, 'h100074, 'h10003c, 'h100075, 'h2004f7, 'h10007a, 'h100077, 'h100047, 'h100078, 'h100079, 'h10007e, 'h10007b, 'h10007c, 'h10007d, 'h100082, 'h10006e, 'h10007f, 'h10006f, 'h100080, 'h100070, 'h100081, 'h100071, 'h100072, 'h10003c, 'h100086, 'h2004f7, 'h100083, 'h100084, 'h100047, 'h100085, 'h10008a, 'h100087, 'h100088, 'h100089, 'h10008e, 'h10008b, 'h10006e, 'h10008c, 'h10006f, 'h10008d, 'h100070, 'h100092, 'h10008f, 'h100090, 'h10003c, 'h100091, 'h2004f7, 'h100071, 'h100072, 'h100047, 'h100096, 'h100093, 'h100094, 'h100095, 'h10009a, 'h100097, 'h100098, 'h100099, 'h10009e, 'h10006e, 'h10009b, 'h10006f, 'h10009c, 'h100070, 'h10009d, 'h10003c, 'h1000a2, 'h2004f7, 'h10009f, 'h1000a0, 'h100047, 'h1000a1, 'h100071, 'h100072, 'h1000a6, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a7, 'h1000aa, 'h10006e, 'h1000a8, 'h10006f, 'h1000a9, 'h100070, 'h1000ab, 'h1000ae, 'h10003c, 'h2004f7, 'h1000ac, 'h1000ad, 'h100047, 'h1000af, 'h1000b2, 'h100072, 'h1000b0, 'h1000b1, 'h100071, 'h1000b3, 'h1000b6, 'h1000b4, 'h1000b5, 'h1000b7, 'h1000ba, 'h10006e, 'h10006f, 'h1000b8, 'h100070, 'h10003c, 'h2004f7, 'h1000b9, 'h1000bb, 'h100047, 'h1000be, 'h1000bc, 'h1000bd, 'h100072, 'h1000bf, 'h1000c2, 'h1000c0, 'h1000c1, 'h100071, 'h1000c3, 'h1000c6, 'h1000c4, 'h1000c5, 'h1000c7, 'h1000ca, 'h10006e, 'h10003c, 'h2004f7, 'h10006f, 'h1000c8, 'h100047, 'h100070, 'h1000c9, 'h1000cb, 'h100072, 'h1000ce, 'h1000cc, 'h1000cd, 'h1000cf, 'h1000d2, 'h1000d0, 'h1000d1, 'h100071, 'h1000d3, 'h1000d6, 'h1000d4, 'h1000d5, 'h10003c, 'h2004f7, 'h1000d7, 'h1000da, 'h100047, 'h10006e, 'h10006f, 'h1000d8, 'h100070, 'h1000d9, 'h100072, 'h1000db, 'h1000df, 'h1000dc, 'h1000dd, 'h1000de, 'h100071, 'h1000e3, 'h1000e0, 'h1000e1, 'h1000e2, 'h10003c, 'h2004f7, 'h1000e7, 'h1000e4, 'h100047, 'h1000e5, 'h1000e6, 'h1000eb, 'h10006e, 'h10006f, 'h1000e8, 'h100070, 'h1000e9, 'h1000ea, 'h100072, 'h1000ef, 'h1000ec, 'h1000ed, 'h100071, 'h1000ee, 'h1000f3, 'h10003c, 'h2004f7, 'h1000f0, 'h1000f1, 'h100047, 'h1000f2, 'h1000f7, 'h1000f4, 'h10006e, 'h10006f, 'h1000f5, 'h100070, 'h1000f6, 'h1000fb, 'h100072, 'h1000f8, 'h1000f9, 'h1000fa, 'h100071, 'h1000ff, 'h1000fc, 'h10003c, 'h2004f7, 'h1000fd, 'h1000fe, 'h100047, 'h100103, 'h100100, 'h100101, 'h100102, 'h100107, 'h10006e, 'h100104, 'h10006f, 'h100105, 'h100070, 'h100106, 'h100072, 'h10010b, 'h100108, 'h100109, 'h10010a, 'h10003c, 'h2004f7, 'h100071, 'h10010f, 'h100047, 'h10010c, 'h10010d, 'h10010e, 'h100113, 'h100110, 'h10006e, 'h100111, 'h10006f, 'h100112, 'h100070, 'h100117, 'h100072, 'h100114, 'h100115, 'h100116, 'h10011b, 'h10003c, 'h2004f7, 'h100118, 'h100119, 'h100047, 'h10011a, 'h100071, 'h10011f, 'h10011c, 'h10011d, 'h10011e, 'h100123, 'h10006e, 'h100120, 'h10006f, 'h100121, 'h100070, 'h100122, 'h100072, 'h100127, 'h100124, 'h10003c, 'h2004f7, 'h100125, 'h100126, 'h100047, 'h100128, 'h10012b, 'h100129, 'h10012a, 'h100071, 'h10012c, 'h10012f, 'h10006e, 'h10012d, 'h10006f, 'h10012e, 'h100070, 'h100130, 'h100072, 'h100133, 'h100131, 'h10003c, 'h2004f7, 'h100132, 'h100134, 'h100047, 'h100137, 'h100135, 'h100136, 'h100138, 'h10013b, 'h100139, 'h10013a, 'h100071, 'h10013c, 'h10013f, 'h10006e, 'h10006f, 'h10013d, 'h100070, 'h10013e, 'h100072, 'h10003c, 'h2004f7, 'h100140, 'h100143, 'h100047, 'h100141, 'h100142, 'h100144, 'h100147, 'h100145, 'h100146, 'h100148, 'h10014b, 'h100149, 'h10014a, 'h100071, 'h10014c, 'h10014f, 'h10006e, 'h10006f, 'h10014d, 'h10003c, 'h2004f7, 'h100070, 'h10014e, 'h100047, 'h100072, 'h100150, 'h100153, 'h100151, 'h100152, 'h100154, 'h100157, 'h100155, 'h100156, 'h100158, 'h10015b, 'h100159, 'h10015a, 'h100071, 'h10015c, 'h100160, 'h10003c, 'h2004f7, 'h10006e, 'h10006f, 'h100047, 'h10015d, 'h100070, 'h10015e, 'h10015f, 'h100072, 'h100164, 'h100161, 'h100162, 'h100163, 'h100168, 'h100165, 'h100166, 'h100167, 'h100071, 'h10016c, 'h100169, 'h10003c, 'h2004f7, 'h10016a, 'h10016b, 'h100047, 'h100170, 'h10006e, 'h10006f, 'h10016d, 'h100070, 'h10016e, 'h10016f, 'h100072, 'h100076, 'h100077, 'h100073, 'h100078, 'h100074, 'h100079, 'h100075, 'h10007a, 'h10003c, 'h2004f7, 'h10007b, 'h10007c, 'h100047, 'h10007d, 'h10007e, 'h10007f, 'h100080, 'h100081, 'h100082, 'h100083, 'h100072, 'h100084, 'h100085, 'h100086, 'h100076, 'h100087, 'h100073, 'h100088, 'h100074, 'h10003c, 'h2004f7, 'h100089, 'h100075, 'h100047, 'h10008a, 'h10008b, 'h10008c, 'h10008d, 'h10008e, 'h10008f, 'h100090, 'h100091, 'h100092, 'h100072, 'h100093, 'h100094, 'h100095, 'h100096, 'h100076, 'h100097, 'h10003c, 'h2004f7, 'h100073, 'h100098, 'h100047, 'h100074, 'h100099, 'h100075, 'h10009a, 'h10009b, 'h10009c, 'h10009d, 'h10009e, 'h10009f, 'h100072, 'h1000a0, 'h1000a1, 'h1000a2, 'h1000a3, 'h100076, 'h1000a4, 'h10003c, 'h2004f7, 'h100073, 'h1000a5, 'h100047, 'h100074, 'h1000a6, 'h100075, 'h1000a7, 'h1000a8, 'h1000a9, 'h1000aa, 'h1000ab, 'h1000ac, 'h1000ad, 'h1000ae, 'h1000af, 'h100072, 'h1000b0, 'h1000b1, 'h1000b2, 'h10003c, 'h2004f7, 'h100076, 'h1000b3, 'h100047, 'h100073, 'h1000b4, 'h100074, 'h1000b5, 'h100075, 'h1000b6, 'h1000b7, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h100072, 'h10003c, 'h2004f7, 'h1000c0, 'h1000c1, 'h100047, 'h1000c2, 'h100076, 'h1000c3, 'h100073, 'h1000c4, 'h100074, 'h1000c5, 'h100075, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h10003c, 'h2004f7, 'h1000ce, 'h1000cf, 'h100047, 'h100072, 'h1000d0, 'h1000d1, 'h1000d2, 'h100076, 'h1000d3, 'h100073, 'h1000d4, 'h100074, 'h1000d5, 'h100075, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h10003c, 'h2004f7, 'h1000db, 'h1000dc, 'h100047, 'h1000dd, 'h1000de, 'h1000df, 'h100072, 'h1000e0, 'h1000e1, 'h1000e2, 'h100076, 'h1000e3, 'h100073, 'h1000e4, 'h100074, 'h1000e5, 'h100075, 'h1000e6, 'h1000e7, 'h10003c, 'h2004f7, 'h1000e8, 'h1000e9, 'h100047, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h100072, 'h1000f0, 'h1000f1, 'h1000f2, 'h100076, 'h1000f3, 'h1000f4, 'h100073, 'h1000f5, 'h100074, 'h10003c, 'h2004f7, 'h1000f6, 'h100075, 'h100047, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h100072, 'h1000fd, 'h1000fe, 'h1000ff, 'h100076, 'h100100, 'h100101, 'h100073, 'h100102, 'h100074, 'h10003c, 'h2004f7, 'h100103, 'h100075, 'h100047, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h100072, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100076, 'h100110, 'h100073, 'h10003c, 'h2004f7, 'h100111, 'h100074, 'h100047, 'h100112, 'h100075, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h100072, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h10003c, 'h2004f7, 'h100076, 'h100120, 'h100047, 'h100073, 'h100121, 'h100074, 'h100122, 'h100075, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h100072, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10003c, 'h2004f7, 'h100076, 'h10012d, 'h100047, 'h100073, 'h10012e, 'h100074, 'h10012f, 'h100075, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100072, 'h100139, 'h10003c, 'h2004f7, 'h10013a, 'h10013b, 'h100047, 'h100076, 'h10013c, 'h100073, 'h10013d, 'h100074, 'h10013e, 'h100075, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h10003c, 'h2004f7, 'h100148, 'h100072, 'h100047, 'h100149, 'h10014a, 'h10014b, 'h100076, 'h10014c, 'h100073, 'h10014d, 'h100074, 'h10014e, 'h100075, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h10003c, 'h2004f7, 'h100155, 'h100156, 'h100047, 'h100157, 'h100158, 'h100072, 'h100159, 'h10015a, 'h10015b, 'h100076, 'h10015c, 'h100073, 'h10015d, 'h100074, 'h10015e, 'h100075, 'h10015f, 'h100160, 'h100161, 'h10003c, 'h2004f7, 'h100162, 'h100163, 'h100047, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100072, 'h100169, 'h10016a, 'h10016b, 'h100076, 'h10016c, 'h100073, 'h10016d, 'h100074, 'h10016e, 'h100075, 'h10003c, 'h2004f7, 'h10016f, 'h100170, 'h100047, 'h10007a, 'h10007b, 'h100077, 'h10007c, 'h100078, 'h10007d, 'h100079, 'h10007e, 'h10007f, 'h100076, 'h100080, 'h100081, 'h100082, 'h100083, 'h100084, 'h100085, 'h10003c, 'h2004f7, 'h100086, 'h100087, 'h100047, 'h100088, 'h100089, 'h10008a, 'h10007a, 'h10008b, 'h100077, 'h10008c, 'h100078, 'h10008d, 'h100079, 'h10008e, 'h100076, 'h10008f, 'h100090, 'h100091, 'h100092, 'h10003c, 'h2004f7, 'h100093, 'h100094, 'h100047, 'h100095, 'h100096, 'h100097, 'h100098, 'h100099, 'h10009a, 'h10007a, 'h10009b, 'h100077, 'h10009c, 'h100078, 'h10009d, 'h100079, 'h10009e, 'h10009f, 'h100076, 'h10003c, 'h2004f7, 'h1000a0, 'h1000a1, 'h100047, 'h1000a2, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h1000a7, 'h10007a, 'h1000a8, 'h100077, 'h1000a9, 'h100078, 'h1000aa, 'h100079, 'h1000ab, 'h1000ac, 'h1000ad, 'h10003c, 'h2004f7, 'h1000ae, 'h1000af, 'h100047, 'h100076, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h10007a, 'h1000b7, 'h100077, 'h1000b8, 'h100078, 'h1000b9, 'h100079, 'h1000ba, 'h10003c, 'h2004f7, 'h1000bb, 'h1000bc, 'h100047, 'h1000bd, 'h1000be, 'h1000bf, 'h100076, 'h1000c0, 'h1000c1, 'h1000c2, 'h1000c3, 'h10007a, 'h1000c4, 'h100077, 'h1000c5, 'h100078, 'h1000c6, 'h100079, 'h1000c7, 'h10003c, 'h2004f7, 'h1000c8, 'h1000c9, 'h100047, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h100076, 'h1000d0, 'h1000d1, 'h1000d2, 'h10007a, 'h1000d3, 'h100077, 'h1000d4, 'h100078, 'h1000d5, 'h10003c, 'h2004f7, 'h100079, 'h1000d6, 'h100047, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h1000df, 'h100076, 'h1000e0, 'h1000e1, 'h1000e2, 'h10007a, 'h1000e3, 'h100077, 'h10003c, 'h2004f7, 'h1000e4, 'h100078, 'h100047, 'h1000e5, 'h100079, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h100076, 'h1000f0, 'h1000f1, 'h1000f2, 'h10003c, 'h2004f7, 'h10007a, 'h1000f3, 'h100047, 'h100077, 'h1000f4, 'h100078, 'h1000f5, 'h100079, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h100076, 'h1000fd, 'h1000fe, 'h1000ff, 'h10003c, 'h2004f7, 'h10007a, 'h100100, 'h100047, 'h100077, 'h100101, 'h100078, 'h100102, 'h100079, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h100076, 'h10010c, 'h10003c, 'h2004f7, 'h10010d, 'h10010e, 'h100047, 'h10010f, 'h10007a, 'h100110, 'h100077, 'h100111, 'h100078, 'h100112, 'h100079, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h100076, 'h100119, 'h10003c, 'h2004f7, 'h10011a, 'h10011b, 'h100047, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h10007a, 'h100120, 'h100077, 'h100121, 'h100078, 'h100122, 'h100079, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h10003c, 'h2004f7, 'h100128, 'h100076, 'h100047, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10007a, 'h10012d, 'h100077, 'h10012e, 'h100078, 'h10012f, 'h100079, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h10003c, 'h2004f7, 'h100135, 'h100136, 'h100047, 'h100137, 'h100138, 'h100076, 'h100139, 'h10013a, 'h10013b, 'h10007a, 'h10013c, 'h100077, 'h10013d, 'h100078, 'h10013e, 'h100079, 'h10013f, 'h100140, 'h100141, 'h10003c, 'h2004f7, 'h100142, 'h100143, 'h100047, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100076, 'h100149, 'h10014a, 'h10014b, 'h10007a, 'h10014c, 'h100077, 'h10014d, 'h100078, 'h10014e, 'h100079, 'h10003c, 'h2004f7, 'h10014f, 'h100150, 'h100047, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100076, 'h100159, 'h10015a, 'h10015b, 'h10007a, 'h10015c, 'h100077, 'h10015d, 'h10003c, 'h2004f7, 'h100078, 'h10015e, 'h100047, 'h100079, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100076, 'h100169, 'h10016a, 'h10016b, 'h10007a, 'h10003c, 'h2004f7, 'h10016c, 'h100077, 'h100047, 'h10016d, 'h100078, 'h10016e, 'h100079, 'h10016f, 'h100170, 'h10007e, 'h10007f, 'h10007b, 'h100080, 'h10007c, 'h100081, 'h10007d, 'h100082, 'h100083, 'h10007a, 'h10003c, 'h2004f7, 'h100084, 'h100085, 'h100047, 'h100086, 'h100087, 'h100088, 'h100089, 'h10008a, 'h10008b, 'h10008c, 'h10008d, 'h10008e, 'h10007e, 'h10008f, 'h10007b, 'h100090, 'h10007c, 'h100091, 'h10007d, 'h10003c, 'h2004f7, 'h100092, 'h10007a, 'h100047, 'h100093, 'h100094, 'h100095, 'h100096, 'h100097, 'h100098, 'h100099, 'h10009a, 'h10009b, 'h10007e, 'h10009c, 'h10007b, 'h10009d, 'h10007c, 'h10009e, 'h10007d, 'h10003c, 'h2004f7, 'h10009f, 'h10007a, 'h100047, 'h1000a0, 'h1000a1, 'h1000a2, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h1000a7, 'h1000a8, 'h1000a9, 'h1000aa, 'h10007e, 'h1000ab, 'h10007b, 'h1000ac, 'h10007c, 'h10003c, 'h2004f7, 'h1000ad, 'h10007d, 'h100047, 'h1000ae, 'h1000af, 'h10007a, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h1000b7, 'h10007e, 'h1000b8, 'h10007b, 'h1000b9, 'h10007c, 'h10003c, 'h2004f7, 'h1000ba, 'h10007d, 'h100047, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h10007a, 'h1000c0, 'h1000c1, 'h1000c2, 'h1000c3, 'h1000c4, 'h1000c5, 'h1000c6, 'h10007e, 'h1000c7, 'h10007b, 'h10003c, 'h2004f7, 'h1000c8, 'h10007c, 'h100047, 'h1000c9, 'h10007d, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h10007a, 'h1000d0, 'h1000d1, 'h1000d2, 'h1000d3, 'h10007e, 'h1000d4, 'h10007b, 'h10003c, 'h2004f7, 'h1000d5, 'h10007c, 'h100047, 'h1000d6, 'h10007d, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h1000df, 'h10007a, 'h1000e0, 'h1000e1, 'h1000e2, 'h10007e, 'h10003c, 'h2004f7, 'h1000e3, 'h10007b, 'h100047, 'h1000e4, 'h10007c, 'h1000e5, 'h10007d, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h10007a, 'h1000f0, 'h10003c, 'h2004f7, 'h1000f1, 'h1000f2, 'h100047, 'h10007e, 'h1000f3, 'h10007b, 'h1000f4, 'h10007c, 'h1000f5, 'h10007d, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h10003c, 'h2004f7, 'h1000ff, 'h10007a, 'h100047, 'h100100, 'h100101, 'h10007b, 'h100102, 'h10007c, 'h100103, 'h10007d, 'h10007e, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10003c, 'h2004f7, 'h10010c, 'h10007a, 'h100047, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h10007b, 'h100111, 'h10007c, 'h100112, 'h10007d, 'h100113, 'h10007e, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h10003c, 'h2004f7, 'h100119, 'h10011a, 'h100047, 'h10011b, 'h10011c, 'h10007a, 'h10011d, 'h10007b, 'h10011e, 'h10007c, 'h10011f, 'h10007d, 'h100120, 'h10007e, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h10003c, 'h2004f7, 'h100126, 'h100127, 'h100047, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10007a, 'h10007b, 'h10012d, 'h10007c, 'h10012e, 'h10007d, 'h10012f, 'h10007e, 'h100130, 'h100131, 'h100132, 'h10003c, 'h2004f7, 'h100133, 'h100134, 'h100047, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10007a, 'h10007b, 'h10013d, 'h10007c, 'h10013e, 'h10007d, 'h10013f, 'h10007e, 'h10003c, 'h2004f7, 'h100140, 'h100141, 'h100047, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10007a, 'h10007b, 'h10014d, 'h10007c, 'h10014e, 'h10003c, 'h2004f7, 'h10007d, 'h10014f, 'h100047, 'h10007e, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10007a, 'h10007b, 'h10003c, 'h2004f7, 'h10015d, 'h10007c, 'h100047, 'h10015e, 'h10007d, 'h10015f, 'h10007e, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10003c, 'h2004f7, 'h10016c, 'h10007a, 'h100047, 'h10007b, 'h10016d, 'h10007c, 'h10016e, 'h10007d, 'h10016f, 'h10007e, 'h100170, 'h100082, 'h100083, 'h10007f, 'h100084, 'h100080, 'h100085, 'h100081, 'h100086, 'h10003c, 'h2004f7, 'h100087, 'h100088, 'h100047, 'h100089, 'h10008a, 'h10008b, 'h10008c, 'h10008d, 'h10008e, 'h10007e, 'h10008f, 'h100090, 'h100091, 'h100092, 'h100082, 'h100093, 'h10007f, 'h100094, 'h100080, 'h10003c, 'h2004f7, 'h100095, 'h100081, 'h100047, 'h100096, 'h100097, 'h100098, 'h100099, 'h10009a, 'h10009b, 'h10007e, 'h10009c, 'h10009d, 'h10009e, 'h10009f, 'h100082, 'h1000a0, 'h10007f, 'h1000a1, 'h100080, 'h10003c, 'h2004f7, 'h1000a2, 'h100081, 'h100047, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h1000a7, 'h1000a8, 'h1000a9, 'h1000aa, 'h1000ab, 'h10007e, 'h1000ac, 'h1000ad, 'h1000ae, 'h100082, 'h1000af, 'h10007f, 'h10003c, 'h2004f7, 'h1000b0, 'h100080, 'h100047, 'h1000b1, 'h100081, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h1000b7, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h10007e, 'h1000bc, 'h1000bd, 'h1000be, 'h10003c, 'h2004f7, 'h100082, 'h1000bf, 'h100047, 'h10007f, 'h1000c0, 'h100080, 'h1000c1, 'h100081, 'h1000c2, 'h1000c3, 'h1000c4, 'h1000c5, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h10007e, 'h10003c, 'h2004f7, 'h1000cc, 'h1000cd, 'h100047, 'h1000ce, 'h100082, 'h1000cf, 'h10007f, 'h1000d0, 'h100080, 'h1000d1, 'h100081, 'h1000d2, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h10003c, 'h2004f7, 'h1000da, 'h1000db, 'h100047, 'h10007e, 'h1000dc, 'h1000dd, 'h1000de, 'h100082, 'h1000df, 'h10007f, 'h1000e0, 'h100080, 'h1000e1, 'h100081, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h10003c, 'h2004f7, 'h1000e7, 'h1000e8, 'h100047, 'h1000e9, 'h1000ea, 'h1000eb, 'h10007e, 'h1000ec, 'h1000ed, 'h1000ee, 'h100082, 'h1000ef, 'h10007f, 'h1000f0, 'h100080, 'h1000f1, 'h100081, 'h1000f2, 'h1000f3, 'h10003c, 'h2004f7, 'h1000f4, 'h1000f5, 'h100047, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h10007e, 'h1000fc, 'h1000fd, 'h1000fe, 'h100082, 'h1000ff, 'h100100, 'h10007f, 'h100101, 'h100080, 'h10003c, 'h2004f7, 'h100102, 'h100081, 'h100047, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h10007e, 'h100109, 'h10010a, 'h10010b, 'h100082, 'h10010c, 'h10010d, 'h10007f, 'h10010e, 'h100080, 'h10003c, 'h2004f7, 'h10010f, 'h100081, 'h100047, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h10007e, 'h100119, 'h10011a, 'h10011b, 'h100082, 'h10011c, 'h10007f, 'h10003c, 'h2004f7, 'h10011d, 'h100080, 'h100047, 'h10011e, 'h100081, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h10007e, 'h100129, 'h10012a, 'h10012b, 'h10003c, 'h2004f7, 'h100082, 'h10012c, 'h100047, 'h10007f, 'h10012d, 'h100080, 'h10012e, 'h100081, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h10007e, 'h10003c, 'h2004f7, 'h100139, 'h10013a, 'h100047, 'h10013b, 'h100082, 'h10013c, 'h10007f, 'h10013d, 'h100080, 'h10013e, 'h100081, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h10003c, 'h2004f7, 'h100147, 'h100148, 'h100047, 'h10007e, 'h100149, 'h10014a, 'h10014b, 'h100082, 'h10014c, 'h10007f, 'h10014d, 'h100080, 'h10014e, 'h100081, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h10003c, 'h2004f7, 'h100154, 'h100155, 'h100047, 'h100156, 'h100157, 'h100158, 'h10007e, 'h100159, 'h10015a, 'h10015b, 'h100082, 'h10015c, 'h10007f, 'h10015d, 'h100080, 'h10015e, 'h100081, 'h10015f, 'h100160, 'h10003c, 'h2004f7, 'h100161, 'h100162, 'h100047, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h10007e, 'h100169, 'h10016a, 'h10016b, 'h100082, 'h10016c, 'h10007f, 'h10016d, 'h100080, 'h10016e, 'h10003c, 'h2004f7, 'h100081, 'h10016f, 'h100047, 'h100170, 'h100086, 'h100087, 'h100083, 'h100088, 'h100084, 'h100089, 'h100085, 'h10008a, 'h10008b, 'h100082, 'h10008c, 'h10008d, 'h10008e, 'h10008f, 'h100090, 'h10003c, 'h2004f7, 'h100091, 'h100092, 'h100047, 'h100093, 'h100086, 'h100094, 'h100083, 'h100095, 'h100084, 'h100096, 'h100085, 'h100097, 'h100098, 'h100099, 'h10009a, 'h10009b, 'h100082, 'h10009c, 'h10009d, 'h10003c, 'h2004f7, 'h10009e, 'h10009f, 'h100047, 'h1000a0, 'h1000a1, 'h1000a2, 'h100086, 'h1000a3, 'h100083, 'h1000a4, 'h100084, 'h1000a5, 'h100085, 'h1000a6, 'h1000a7, 'h1000a8, 'h1000a9, 'h1000aa, 'h1000ab, 'h10003c, 'h2004f7, 'h100082, 'h1000ac, 'h100047, 'h1000ad, 'h1000ae, 'h1000af, 'h100086, 'h1000b0, 'h100083, 'h1000b1, 'h100084, 'h1000b2, 'h100085, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h1000b7, 'h1000b8, 'h10003c, 'h2004f7, 'h1000b9, 'h1000ba, 'h100047, 'h1000bb, 'h100082, 'h1000bc, 'h1000bd, 'h1000be, 'h100086, 'h1000bf, 'h100083, 'h1000c0, 'h100084, 'h1000c1, 'h100085, 'h1000c2, 'h1000c3, 'h1000c4, 'h1000c5, 'h10003c, 'h2004f7, 'h1000c6, 'h1000c7, 'h100047, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h100082, 'h1000cc, 'h1000cd, 'h1000ce, 'h100086, 'h1000cf, 'h100083, 'h1000d0, 'h100084, 'h1000d1, 'h100085, 'h1000d2, 'h10003c, 'h2004f7, 'h1000d3, 'h1000d4, 'h100047, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h100082, 'h1000dc, 'h1000dd, 'h1000de, 'h100086, 'h1000df, 'h100083, 'h1000e0, 'h100084, 'h10003c, 'h2004f7, 'h1000e1, 'h100085, 'h100047, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h100082, 'h1000ec, 'h1000ed, 'h1000ee, 'h100086, 'h1000ef, 'h10003c, 'h2004f7, 'h100083, 'h1000f0, 'h100047, 'h100084, 'h1000f1, 'h100085, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h100082, 'h1000fc, 'h1000fd, 'h10003c, 'h2004f7, 'h1000fe, 'h100086, 'h100047, 'h1000ff, 'h100083, 'h100100, 'h100084, 'h100101, 'h100085, 'h100102, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100082, 'h100109, 'h10010a, 'h10003c, 'h2004f7, 'h10010b, 'h100086, 'h100047, 'h10010c, 'h100083, 'h10010d, 'h100084, 'h10010e, 'h100085, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h10003c, 'h2004f7, 'h100082, 'h100119, 'h100047, 'h10011a, 'h10011b, 'h100086, 'h10011c, 'h100083, 'h10011d, 'h100084, 'h10011e, 'h100085, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h10003c, 'h2004f7, 'h100126, 'h100127, 'h100047, 'h100128, 'h100082, 'h100129, 'h10012a, 'h10012b, 'h100086, 'h10012c, 'h100083, 'h10012d, 'h100084, 'h10012e, 'h100085, 'h10012f, 'h100130, 'h100131, 'h100132, 'h10003c, 'h2004f7, 'h100133, 'h100134, 'h100047, 'h100135, 'h100136, 'h100137, 'h100138, 'h100082, 'h100139, 'h10013a, 'h10013b, 'h100086, 'h10013c, 'h100083, 'h10013d, 'h100084, 'h10013e, 'h100085, 'h10013f, 'h10003c, 'h2004f7, 'h100140, 'h100141, 'h100047, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100082, 'h100149, 'h10014a, 'h10014b, 'h100086, 'h10014c, 'h100083, 'h10014d, 'h100084, 'h10003c, 'h2004f7, 'h10014e, 'h100085, 'h100047, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100082, 'h100159, 'h10015a, 'h10015b, 'h100086, 'h10015c, 'h10003c, 'h2004f7, 'h100083, 'h10015d, 'h100047, 'h100084, 'h10015e, 'h100085, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100082, 'h100169, 'h10016a, 'h10003c, 'h2004f7, 'h10016b, 'h100086, 'h100047, 'h10016c, 'h100083, 'h10016d, 'h100084, 'h10016e, 'h100085, 'h10016f, 'h100170, 'h10008a, 'h10008b, 'h100087, 'h10008c, 'h100088, 'h10008d, 'h100089, 'h10008e, 'h10003c, 'h2004f7, 'h10008f, 'h100086, 'h100047, 'h100090, 'h100091, 'h100092, 'h100093, 'h100094, 'h100095, 'h100096, 'h100097, 'h10008a, 'h100098, 'h100087, 'h100099, 'h100088, 'h10009a, 'h100089, 'h10009b, 'h10003c, 'h2004f7, 'h10009c, 'h10009d, 'h100047, 'h10009e, 'h10009f, 'h100086, 'h1000a0, 'h1000a1, 'h1000a2, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h10008a, 'h1000a7, 'h100087, 'h1000a8, 'h100088, 'h1000a9, 'h10003c, 'h2004f7, 'h100089, 'h1000aa, 'h100047, 'h1000ab, 'h1000ac, 'h1000ad, 'h1000ae, 'h1000af, 'h100086, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h10008a, 'h1000b4, 'h100087, 'h1000b5, 'h100088, 'h1000b6, 'h10003c, 'h2004f7, 'h100089, 'h1000b7, 'h100047, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h100086, 'h1000c0, 'h1000c1, 'h1000c2, 'h10008a, 'h1000c3, 'h100087, 'h1000c4, 'h10003c, 'h2004f7, 'h100088, 'h1000c5, 'h100047, 'h100089, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h100086, 'h1000d0, 'h1000d1, 'h1000d2, 'h10008a, 'h10003c, 'h2004f7, 'h1000d3, 'h100087, 'h100047, 'h1000d4, 'h100088, 'h1000d5, 'h100089, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h1000df, 'h100086, 'h1000e0, 'h10003c, 'h2004f7, 'h1000e1, 'h1000e2, 'h100047, 'h10008a, 'h1000e3, 'h100087, 'h1000e4, 'h100088, 'h1000e5, 'h100089, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h10003c, 'h2004f7, 'h1000ef, 'h100086, 'h100047, 'h1000f0, 'h1000f1, 'h1000f2, 'h10008a, 'h1000f3, 'h100087, 'h1000f4, 'h100088, 'h1000f5, 'h100089, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h10003c, 'h2004f7, 'h1000fc, 'h1000fd, 'h100047, 'h1000fe, 'h1000ff, 'h100086, 'h100100, 'h100101, 'h100102, 'h10008a, 'h100103, 'h100087, 'h100104, 'h100088, 'h100105, 'h100089, 'h100106, 'h100107, 'h100108, 'h10003c, 'h2004f7, 'h100109, 'h10010a, 'h100047, 'h10010b, 'h10010c, 'h100086, 'h10010d, 'h10010e, 'h10010f, 'h10008a, 'h100110, 'h100087, 'h100111, 'h100088, 'h100112, 'h100089, 'h100113, 'h100114, 'h100115, 'h10003c, 'h2004f7, 'h100116, 'h100117, 'h100047, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h100086, 'h10011d, 'h10011e, 'h10011f, 'h10008a, 'h100120, 'h100087, 'h100121, 'h100088, 'h100122, 'h100089, 'h10003c, 'h2004f7, 'h100123, 'h100124, 'h100047, 'h100125, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h100086, 'h10012d, 'h10012e, 'h10012f, 'h10008a, 'h100130, 'h100087, 'h100131, 'h10003c, 'h2004f7, 'h100088, 'h100132, 'h100047, 'h100089, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h100086, 'h10013d, 'h10013e, 'h10013f, 'h10008a, 'h10003c, 'h2004f7, 'h100140, 'h100087, 'h100047, 'h100141, 'h100088, 'h100142, 'h100089, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h100086, 'h10014d, 'h10003c, 'h2004f7, 'h10014e, 'h10014f, 'h100047, 'h10008a, 'h100150, 'h100087, 'h100151, 'h100088, 'h100152, 'h100089, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10003c, 'h2004f7, 'h10015c, 'h100086, 'h100047, 'h10015d, 'h10015e, 'h10015f, 'h10008a, 'h100160, 'h100087, 'h100161, 'h100088, 'h100162, 'h100089, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h10003c, 'h2004f7, 'h100169, 'h10016a, 'h100047, 'h10016b, 'h10016c, 'h100086, 'h10016d, 'h10016e, 'h10016f, 'h10008a, 'h100170, 'h10008f, 'h10008e, 'h10008b, 'h100090, 'h10008c, 'h100091, 'h10008d, 'h100092, 'h10003c, 'h2004f7, 'h100093, 'h100094, 'h100047, 'h100095, 'h100096, 'h100097, 'h100098, 'h100099, 'h10009a, 'h10009b, 'h10009c, 'h10009d, 'h10009e, 'h10008e, 'h10009f, 'h10008b, 'h1000a0, 'h10008c, 'h1000a1, 'h10003c, 'h2004f7, 'h10008d, 'h1000a2, 'h100047, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h1000a7, 'h1000a8, 'h1000a9, 'h1000aa, 'h1000ab, 'h1000ac, 'h1000ad, 'h1000ae, 'h10008e, 'h1000af, 'h10008b, 'h1000b0, 'h10003c, 'h2004f7, 'h10008c, 'h1000b1, 'h100047, 'h10008d, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h1000b7, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h10008e, 'h1000bf, 'h10003c, 'h2004f7, 'h10008b, 'h1000c0, 'h100047, 'h10008c, 'h1000c1, 'h10008d, 'h1000c2, 'h1000c3, 'h1000c4, 'h1000c5, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h10003c, 'h2004f7, 'h10008e, 'h1000cf, 'h100047, 'h10008b, 'h1000d0, 'h10008c, 'h1000d1, 'h10008d, 'h1000d2, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h10003c, 'h2004f7, 'h1000dd, 'h1000de, 'h100047, 'h10008e, 'h1000df, 'h10008b, 'h1000e0, 'h10008c, 'h1000e1, 'h10008d, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h10003c, 'h2004f7, 'h1000eb, 'h1000ec, 'h100047, 'h1000ed, 'h1000ee, 'h10008e, 'h1000ef, 'h10008b, 'h1000f0, 'h10008c, 'h1000f1, 'h10008d, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h10003c, 'h2004f7, 'h1000f9, 'h1000fa, 'h100047, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h10008e, 'h1000ff, 'h10008b, 'h100100, 'h10008c, 'h100101, 'h10008d, 'h100102, 'h100103, 'h100104, 'h100105, 'h100106, 'h10003c, 'h2004f7, 'h100107, 'h100108, 'h100047, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h10008e, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h10008b, 'h100111, 'h10008c, 'h100112, 'h10008d, 'h100113, 'h100114, 'h10003c, 'h2004f7, 'h100115, 'h100116, 'h100047, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10008e, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h10008b, 'h100121, 'h10008c, 'h100122, 'h10008d, 'h10003c, 'h2004f7, 'h100123, 'h100124, 'h100047, 'h100125, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10008e, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h10008b, 'h100131, 'h10008c, 'h10003c, 'h2004f7, 'h100132, 'h10008d, 'h100047, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10008e, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h10008b, 'h10003c, 'h2004f7, 'h100141, 'h10008c, 'h100047, 'h100142, 'h10008d, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10008e, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h10003c, 'h2004f7, 'h100150, 'h10008b, 'h100047, 'h100151, 'h10008c, 'h100152, 'h10008d, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10008e, 'h10015c, 'h10015d, 'h10003c, 'h2004f7, 'h10015e, 'h10015f, 'h100047, 'h100160, 'h10008b, 'h100161, 'h10008c, 'h100162, 'h10008d, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10008e, 'h10003c, 'h2004f7, 'h10016c, 'h10016d, 'h100047, 'h10016e, 'h10016f, 'h100170, 'h100093, 'h100092, 'h10008f, 'h100094, 'h100090, 'h100095, 'h100091, 'h100096, 'h100097, 'h100098, 'h100099, 'h10009a, 'h10009b, 'h10003c, 'h2004f7, 'h10009c, 'h10009d, 'h100047, 'h10009e, 'h10009f, 'h1000a0, 'h1000a1, 'h1000a2, 'h100092, 'h1000a3, 'h10008f, 'h1000a4, 'h100090, 'h1000a5, 'h100091, 'h1000a6, 'h1000a7, 'h1000a8, 'h1000a9, 'h10003c, 'h2004f7, 'h1000aa, 'h1000ab, 'h100047, 'h1000ac, 'h1000ad, 'h1000ae, 'h1000af, 'h1000b0, 'h1000b1, 'h1000b2, 'h100092, 'h1000b3, 'h10008f, 'h1000b4, 'h100090, 'h1000b5, 'h100091, 'h1000b6, 'h1000b7, 'h10003c, 'h2004f7, 'h1000b8, 'h1000b9, 'h100047, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h1000c0, 'h1000c1, 'h1000c2, 'h100092, 'h1000c3, 'h10008f, 'h1000c4, 'h100090, 'h1000c5, 'h100091, 'h10003c, 'h2004f7, 'h1000c6, 'h1000c7, 'h100047, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h1000d0, 'h1000d1, 'h1000d2, 'h100092, 'h1000d3, 'h10008f, 'h1000d4, 'h100090, 'h10003c, 'h2004f7, 'h1000d5, 'h100091, 'h100047, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h1000df, 'h1000e0, 'h1000e1, 'h1000e2, 'h100092, 'h1000e3, 'h10008f, 'h10003c, 'h2004f7, 'h1000e4, 'h100090, 'h100047, 'h1000e5, 'h100091, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h100092, 'h10003c, 'h2004f7, 'h1000f3, 'h10008f, 'h100047, 'h1000f4, 'h100090, 'h1000f5, 'h100091, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h10003c, 'h2004f7, 'h100102, 'h100092, 'h100047, 'h100103, 'h100104, 'h10008f, 'h100090, 'h100105, 'h100091, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h10003c, 'h2004f7, 'h100110, 'h100092, 'h100047, 'h100111, 'h100112, 'h100113, 'h100114, 'h10008f, 'h100115, 'h100090, 'h100116, 'h100091, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10003c, 'h2004f7, 'h10011e, 'h10011f, 'h100047, 'h100092, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h10008f, 'h100125, 'h100090, 'h100126, 'h100091, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10003c, 'h2004f7, 'h10012c, 'h10012d, 'h100047, 'h10012e, 'h10012f, 'h100092, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h10008f, 'h100135, 'h100090, 'h100136, 'h100091, 'h100137, 'h100138, 'h100139, 'h10003c, 'h2004f7, 'h10013a, 'h10013b, 'h100047, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100092, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h10008f, 'h100145, 'h100090, 'h100146, 'h100091, 'h100147, 'h10003c, 'h2004f7, 'h100148, 'h100149, 'h100047, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100092, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h10008f, 'h100155, 'h100090, 'h100156, 'h10003c, 'h2004f7, 'h100091, 'h100157, 'h100047, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100092, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h10008f, 'h100165, 'h10003c, 'h2004f7, 'h100090, 'h100166, 'h100047, 'h100091, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100092, 'h100170, 'h100097, 'h100096, 'h100093, 'h100098, 'h10003c, 'h2004f7, 'h100094, 'h100099, 'h100047, 'h100095, 'h10009a, 'h10009b, 'h10009c, 'h10009d, 'h10009e, 'h10009f, 'h1000a0, 'h1000a1, 'h1000a2, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h100096, 'h1000a7, 'h10003c, 'h2004f7, 'h100093, 'h1000a8, 'h100047, 'h100094, 'h1000a9, 'h100095, 'h1000aa, 'h1000ab, 'h1000ac, 'h1000ad, 'h1000ae, 'h1000af, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h10003c, 'h2004f7, 'h100096, 'h1000b7, 'h100047, 'h100093, 'h1000b8, 'h100094, 'h1000b9, 'h100095, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h1000c0, 'h1000c1, 'h1000c2, 'h1000c3, 'h1000c4, 'h10003c, 'h2004f7, 'h1000c5, 'h1000c6, 'h100047, 'h100096, 'h1000c7, 'h100093, 'h1000c8, 'h100094, 'h1000c9, 'h100095, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h1000d0, 'h1000d1, 'h1000d2, 'h10003c, 'h2004f7, 'h1000d3, 'h1000d4, 'h100047, 'h1000d5, 'h1000d6, 'h100096, 'h1000d7, 'h100093, 'h1000d8, 'h100094, 'h1000d9, 'h100095, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h1000df, 'h1000e0, 'h10003c, 'h2004f7, 'h1000e1, 'h1000e2, 'h100047, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h100096, 'h1000e7, 'h100093, 'h1000e8, 'h100094, 'h1000e9, 'h100095, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h10003c, 'h2004f7, 'h1000ef, 'h1000f0, 'h100047, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h100096, 'h1000f7, 'h100093, 'h1000f8, 'h100094, 'h1000f9, 'h100095, 'h1000fa, 'h1000fb, 'h1000fc, 'h10003c, 'h2004f7, 'h1000fd, 'h1000fe, 'h100047, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100096, 'h100105, 'h100106, 'h100107, 'h100108, 'h100093, 'h100094, 'h100109, 'h100095, 'h10010a, 'h10003c, 'h2004f7, 'h10010b, 'h10010c, 'h100047, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100096, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h100093, 'h100119, 'h100094, 'h10003c, 'h2004f7, 'h10011a, 'h100095, 'h100047, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100096, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h100093, 'h10003c, 'h2004f7, 'h100129, 'h100094, 'h100047, 'h10012a, 'h100095, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100096, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h10003c, 'h2004f7, 'h100138, 'h100093, 'h100047, 'h100139, 'h100094, 'h10013a, 'h100095, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100096, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h10003c, 'h2004f7, 'h100146, 'h100147, 'h100047, 'h100148, 'h100093, 'h100149, 'h100094, 'h10014a, 'h100095, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100096, 'h100150, 'h100151, 'h100152, 'h100153, 'h10003c, 'h2004f7, 'h100154, 'h100155, 'h100047, 'h100156, 'h100157, 'h100158, 'h100093, 'h100159, 'h100094, 'h10015a, 'h100095, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100096, 'h100160, 'h100161, 'h10003c, 'h2004f7, 'h100162, 'h100163, 'h100047, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100093, 'h100169, 'h100094, 'h10016a, 'h100095, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100096, 'h10003c, 'h2004f7, 'h100170, 'h10009b, 'h10009a, 'h100047, 'h100097, 'h10009c, 'h100098, 'h10009d, 'h100099, 'h10009e, 'h10009f, 'h1000a0, 'h1000a1, 'h1000a2, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h1000a7, 'h10003c, 'h2004f7, 'h1000a8, 'h1000a9, 'h1000aa, 'h100047, 'h10009a, 'h1000ab, 'h100097, 'h1000ac, 'h100098, 'h1000ad, 'h100099, 'h1000ae, 'h1000af, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h10003c, 'h2004f7, 'h1000b6, 'h1000b7, 'h1000b8, 'h100047, 'h1000b9, 'h1000ba, 'h10009a, 'h1000bb, 'h100097, 'h1000bc, 'h100098, 'h1000bd, 'h100099, 'h1000be, 'h1000bf, 'h1000c0, 'h1000c1, 'h1000c2, 'h1000c3, 'h10003c, 'h2004f7, 'h1000c4, 'h1000c5, 'h1000c6, 'h100047, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h10009a, 'h1000cb, 'h100097, 'h1000cc, 'h100098, 'h1000cd, 'h100099, 'h1000ce, 'h1000cf, 'h1000d0, 'h1000d1, 'h10003c, 'h2004f7, 'h1000d2, 'h1000d3, 'h1000d4, 'h100047, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h10009a, 'h1000db, 'h100097, 'h1000dc, 'h100098, 'h1000dd, 'h100099, 'h1000de, 'h1000df, 'h10003c, 'h2004f7, 'h1000e0, 'h1000e1, 'h1000e2, 'h100047, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h10009a, 'h1000eb, 'h100097, 'h1000ec, 'h100098, 'h1000ed, 'h100099, 'h10003c, 'h2004f7, 'h1000ee, 'h1000ef, 'h1000f0, 'h100047, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h10009a, 'h1000fb, 'h1000fc, 'h100097, 'h100098, 'h10003c, 'h2004f7, 'h1000fd, 'h100099, 'h1000fe, 'h100047, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h10009a, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h10003c, 'h2004f7, 'h100097, 'h100098, 'h10010d, 'h100047, 'h100099, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h10009a, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10003c, 'h2004f7, 'h10011b, 'h10011c, 'h100097, 'h100047, 'h10011d, 'h100098, 'h10011e, 'h100099, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h10009a, 'h100125, 'h100126, 'h100127, 'h100128, 'h10003c, 'h2004f7, 'h100129, 'h10012a, 'h10012b, 'h100047, 'h10012c, 'h100097, 'h10012d, 'h100098, 'h10012e, 'h100099, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h10009a, 'h100134, 'h100135, 'h100136, 'h10003c, 'h2004f7, 'h100137, 'h100138, 'h100139, 'h100047, 'h10013a, 'h10013b, 'h10013c, 'h100097, 'h10013d, 'h100098, 'h10013e, 'h100099, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h10009a, 'h100144, 'h10003c, 'h2004f7, 'h100145, 'h100146, 'h100147, 'h100047, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h100097, 'h10014d, 'h100098, 'h10014e, 'h100099, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h10003c, 'h2004f7, 'h10009a, 'h100154, 'h100155, 'h100047, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h100097, 'h10015d, 'h100098, 'h10015e, 'h100099, 'h10015f, 'h100160, 'h100161, 'h10003c, 'h2004f7, 'h100162, 'h100163, 'h10009a, 'h100047, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h100097, 'h10016d, 'h100098, 'h10016e, 'h100099, 'h10016f, 'h10003c, 'h2004f7, 'h100170, 'h10009f, 'h10009e, 'h100047, 'h10009b, 'h1000a0, 'h10009c, 'h1000a1, 'h10009d, 'h1000a2, 'h1000a3, 'h1000a4, 'h1000a5, 'h1000a6, 'h1000a7, 'h1000a8, 'h1000a9, 'h1000aa, 'h1000ab, 'h10003c, 'h2004f7, 'h1000ac, 'h1000ad, 'h1000ae, 'h100047, 'h10009e, 'h1000af, 'h10009b, 'h1000b0, 'h10009c, 'h1000b1, 'h10009d, 'h1000b2, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h1000b7, 'h1000b8, 'h1000b9, 'h10003c, 'h2004f7, 'h1000ba, 'h1000bb, 'h1000bc, 'h100047, 'h1000bd, 'h1000be, 'h10009e, 'h1000bf, 'h10009b, 'h1000c0, 'h10009c, 'h1000c1, 'h10009d, 'h1000c2, 'h1000c3, 'h1000c4, 'h1000c5, 'h1000c6, 'h1000c7, 'h10003c, 'h2004f7, 'h1000c8, 'h1000c9, 'h1000ca, 'h100047, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h10009e, 'h1000cf, 'h10009b, 'h1000d0, 'h10009c, 'h1000d1, 'h10009d, 'h1000d2, 'h1000d3, 'h1000d4, 'h1000d5, 'h10003c, 'h2004f7, 'h1000d6, 'h1000d7, 'h1000d8, 'h100047, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h10009e, 'h1000df, 'h10009b, 'h1000e0, 'h10009c, 'h1000e1, 'h10009d, 'h1000e2, 'h1000e3, 'h10003c, 'h2004f7, 'h1000e4, 'h1000e5, 'h1000e6, 'h100047, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h10009e, 'h1000ef, 'h10009b, 'h1000f0, 'h10009c, 'h1000f1, 'h10009d, 'h10003c, 'h2004f7, 'h1000f2, 'h1000f3, 'h1000f4, 'h100047, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h10009e, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h10009b, 'h10009c, 'h10003c, 'h2004f7, 'h100101, 'h10009d, 'h100102, 'h100047, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10009e, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h10003c, 'h2004f7, 'h10009b, 'h10009c, 'h100111, 'h100047, 'h10009d, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h10009e, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10003c, 'h2004f7, 'h10011f, 'h100120, 'h10009b, 'h100047, 'h100121, 'h10009c, 'h100122, 'h10009d, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h10009e, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10003c, 'h2004f7, 'h10012d, 'h10012e, 'h10012f, 'h100047, 'h100130, 'h10009b, 'h100131, 'h10009c, 'h100132, 'h10009d, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h10009e, 'h100138, 'h100139, 'h10013a, 'h10003c, 'h2004f7, 'h10013b, 'h10013c, 'h10013d, 'h100047, 'h10013e, 'h10013f, 'h100140, 'h10009b, 'h100141, 'h10009c, 'h100142, 'h10009d, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h10009e, 'h100148, 'h10003c, 'h2004f7, 'h100149, 'h10014a, 'h10014b, 'h100047, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h10009b, 'h100151, 'h10009c, 'h100152, 'h10009d, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h10003c, 'h2004f7, 'h10009e, 'h100158, 'h100159, 'h100047, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h10009b, 'h100161, 'h10009c, 'h100162, 'h10009d, 'h100163, 'h100164, 'h100165, 'h10003c, 'h2004f7, 'h100166, 'h100167, 'h10009e, 'h100047, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h1000a3, 'h1000a2, 'h10009f, 'h1000a4, 'h1000a0, 'h1000a5, 'h10003c, 'h2004f7, 'h1000a1, 'h1000a6, 'h1000a7, 'h100047, 'h1000a8, 'h1000a9, 'h1000aa, 'h1000ab, 'h1000ac, 'h1000ad, 'h1000ae, 'h1000af, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000a2, 'h1000b3, 'h10009f, 'h1000b4, 'h10003c, 'h2004f7, 'h1000a0, 'h1000b5, 'h1000a1, 'h100047, 'h1000b6, 'h1000b7, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h1000c0, 'h1000c1, 'h1000c2, 'h1000a2, 'h1000c3, 'h10003c, 'h2004f7, 'h10009f, 'h1000c4, 'h1000a0, 'h100047, 'h1000c5, 'h1000a1, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h1000d0, 'h1000d1, 'h1000d2, 'h10003c, 'h2004f7, 'h1000a2, 'h1000d3, 'h10009f, 'h100047, 'h1000d4, 'h1000a0, 'h1000d5, 'h1000a1, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h1000df, 'h1000e0, 'h10003c, 'h2004f7, 'h1000e1, 'h1000e2, 'h1000a2, 'h100047, 'h1000e3, 'h10009f, 'h1000e4, 'h1000a0, 'h1000e5, 'h1000a1, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h10003c, 'h2004f7, 'h1000ef, 'h1000f0, 'h1000f1, 'h100047, 'h1000f2, 'h1000a2, 'h1000f3, 'h1000f4, 'h10009f, 'h1000a0, 'h1000f5, 'h1000a1, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h10003c, 'h2004f7, 'h1000fd, 'h1000fe, 'h1000ff, 'h100047, 'h100100, 'h1000a2, 'h100101, 'h100102, 'h100103, 'h100104, 'h10009f, 'h1000a0, 'h100105, 'h1000a1, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10003c, 'h2004f7, 'h10010b, 'h10010c, 'h10010d, 'h100047, 'h10010e, 'h1000a2, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h10009f, 'h1000a0, 'h100115, 'h1000a1, 'h100116, 'h100117, 'h100118, 'h10003c, 'h2004f7, 'h100119, 'h10011a, 'h10011b, 'h100047, 'h10011c, 'h1000a2, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h10009f, 'h100125, 'h1000a0, 'h100126, 'h1000a1, 'h10003c, 'h2004f7, 'h100127, 'h100128, 'h100129, 'h100047, 'h10012a, 'h10012b, 'h1000a2, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h10009f, 'h100135, 'h1000a0, 'h10003c, 'h2004f7, 'h100136, 'h1000a1, 'h100137, 'h100047, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h1000a2, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h10009f, 'h10003c, 'h2004f7, 'h100145, 'h1000a0, 'h100146, 'h100047, 'h1000a1, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h1000a2, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h10003c, 'h2004f7, 'h100154, 'h10009f, 'h100155, 'h100047, 'h1000a0, 'h100156, 'h1000a1, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h1000a2, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h10003c, 'h2004f7, 'h100162, 'h100163, 'h100164, 'h100047, 'h10009f, 'h100165, 'h1000a0, 'h100166, 'h1000a1, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h1000a2, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h10003c, 'h2004f7, 'h100170, 'h1000a7, 'h1000a6, 'h100047, 'h1000a3, 'h1000a8, 'h1000a4, 'h1000a9, 'h1000a5, 'h1000aa, 'h1000ab, 'h1000ac, 'h1000ad, 'h1000ae, 'h1000af, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h10003c, 'h2004f7, 'h1000b4, 'h1000b5, 'h1000b6, 'h100047, 'h1000a6, 'h1000b7, 'h1000a3, 'h1000b8, 'h1000a4, 'h1000b9, 'h1000a5, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h1000c0, 'h1000c1, 'h10003c, 'h2004f7, 'h1000c2, 'h1000c3, 'h1000c4, 'h100047, 'h1000c5, 'h1000c6, 'h1000a6, 'h1000c7, 'h1000a3, 'h1000c8, 'h1000a4, 'h1000c9, 'h1000a5, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h10003c, 'h2004f7, 'h1000d0, 'h1000d1, 'h1000d2, 'h100047, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000a6, 'h1000d7, 'h1000a3, 'h1000d8, 'h1000a4, 'h1000d9, 'h1000a5, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h10003c, 'h2004f7, 'h1000de, 'h1000df, 'h1000e0, 'h100047, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000a6, 'h1000e7, 'h1000a3, 'h1000e8, 'h1000a4, 'h1000e9, 'h1000a5, 'h1000ea, 'h1000eb, 'h10003c, 'h2004f7, 'h1000ec, 'h1000ed, 'h1000ee, 'h100047, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000a6, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000a3, 'h1000a4, 'h1000f9, 'h1000a5, 'h10003c, 'h2004f7, 'h1000fa, 'h1000fb, 'h1000fc, 'h100047, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h1000a6, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h1000a3, 'h1000a4, 'h10003c, 'h2004f7, 'h100109, 'h1000a5, 'h10010a, 'h100047, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h1000a6, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h10003c, 'h2004f7, 'h1000a3, 'h1000a4, 'h100119, 'h100047, 'h1000a5, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h1000a6, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h100126, 'h10003c, 'h2004f7, 'h100127, 'h100128, 'h1000a3, 'h100047, 'h100129, 'h1000a4, 'h10012a, 'h1000a5, 'h10012b, 'h10012c, 'h1000a6, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h10003c, 'h2004f7, 'h100135, 'h100136, 'h100137, 'h100047, 'h100138, 'h1000a3, 'h100139, 'h1000a4, 'h10013a, 'h1000a5, 'h10013b, 'h1000a6, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h10003c, 'h2004f7, 'h100143, 'h100144, 'h100145, 'h100047, 'h100146, 'h100147, 'h100148, 'h1000a3, 'h100149, 'h1000a4, 'h10014a, 'h1000a5, 'h10014b, 'h1000a6, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h10003c, 'h2004f7, 'h100151, 'h100152, 'h100153, 'h100047, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h1000a3, 'h100159, 'h1000a4, 'h10015a, 'h1000a5, 'h10015b, 'h1000a6, 'h10015c, 'h10015d, 'h10015e, 'h10003c, 'h2004f7, 'h10015f, 'h100160, 'h100161, 'h100047, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h1000a3, 'h100169, 'h1000a4, 'h10016a, 'h1000a5, 'h10016b, 'h1000a6, 'h10016c, 'h10003c, 'h2004f7, 'h10016d, 'h10016e, 'h10016f, 'h100047, 'h100170, 'h1000ab, 'h1000a7, 'h1000ac, 'h1000a8, 'h1000ad, 'h1000a9, 'h1000ae, 'h1000aa, 'h1000af, 'h1000b0, 'h1000b1, 'h1000b2, 'h1000b3, 'h1000b4, 'h10003c, 'h2004f7, 'h1000b5, 'h1000b6, 'h1000b7, 'h100047, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h1000ab, 'h1000a7, 'h1000bc, 'h1000a8, 'h1000bd, 'h1000a9, 'h1000be, 'h1000aa, 'h1000bf, 'h1000c0, 'h1000c1, 'h10003c, 'h2004f7, 'h1000c2, 'h1000c3, 'h1000c4, 'h100047, 'h1000c5, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000ab, 'h1000a7, 'h1000cc, 'h1000a8, 'h1000cd, 'h1000a9, 'h1000ce, 'h1000aa, 'h10003c, 'h2004f7, 'h1000cf, 'h1000d0, 'h1000d1, 'h100047, 'h1000d2, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000ab, 'h1000a7, 'h1000d9, 'h1000a8, 'h1000da, 'h1000a9, 'h1000db, 'h1000aa, 'h10003c, 'h2004f7, 'h1000dc, 'h1000dd, 'h1000de, 'h100047, 'h1000df, 'h1000e0, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000ab, 'h1000e8, 'h1000a7, 'h1000a8, 'h1000e9, 'h1000a9, 'h10003c, 'h2004f7, 'h1000ea, 'h1000aa, 'h1000eb, 'h100047, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000ab, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000a7, 'h10003c, 'h2004f7, 'h1000a8, 'h1000f9, 'h1000a9, 'h100047, 'h1000fa, 'h1000aa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h1000ab, 'h100105, 'h100106, 'h10003c, 'h2004f7, 'h100107, 'h100108, 'h1000a7, 'h100047, 'h1000a8, 'h100109, 'h1000a9, 'h10010a, 'h1000aa, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h1000ab, 'h10003c, 'h2004f7, 'h100115, 'h100116, 'h100047, 'h100117, 'h100118, 'h1000a7, 'h1000a8, 'h100119, 'h1000a9, 'h10011a, 'h1000aa, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h10003c, 'h2004f7, 'h100123, 'h100124, 'h1000ab, 'h100047, 'h100125, 'h100126, 'h100127, 'h100128, 'h1000a7, 'h100129, 'h1000a8, 'h10012a, 'h1000a9, 'h10012b, 'h1000aa, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h10003c, 'h2004f7, 'h100130, 'h100131, 'h100132, 'h100047, 'h100133, 'h100134, 'h1000ab, 'h100135, 'h1000a7, 'h100136, 'h1000a8, 'h100137, 'h1000a9, 'h100138, 'h1000aa, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10003c, 'h2004f7, 'h10013d, 'h10013e, 'h10013f, 'h100047, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h1000ab, 'h1000a7, 'h100145, 'h1000a8, 'h100146, 'h1000a9, 'h100147, 'h1000aa, 'h100148, 'h100149, 'h10003c, 'h2004f7, 'h10014a, 'h10014b, 'h10014c, 'h100047, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h1000ab, 'h1000a7, 'h100155, 'h1000a8, 'h100156, 'h1000a9, 'h100157, 'h10003c, 'h2004f7, 'h1000aa, 'h100158, 'h100159, 'h100047, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h1000ab, 'h1000a7, 'h100162, 'h1000a8, 'h100163, 'h1000a9, 'h100164, 'h10003c, 'h2004f7, 'h1000aa, 'h100165, 'h100166, 'h100047, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h1000af, 'h1000ab, 'h1000b0, 'h1000ac, 'h1000b1, 'h10003c, 'h2004f7, 'h1000ad, 'h1000b2, 'h1000ae, 'h100047, 'h1000b3, 'h1000b4, 'h1000b5, 'h1000b6, 'h1000b7, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h1000af, 'h1000ab, 'h10003c, 'h2004f7, 'h1000c0, 'h1000ac, 'h1000c1, 'h100047, 'h1000ad, 'h1000c2, 'h1000ae, 'h1000c3, 'h1000c4, 'h1000c5, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h10003c, 'h2004f7, 'h1000cf, 'h1000af, 'h1000ab, 'h100047, 'h1000d0, 'h1000ac, 'h1000d1, 'h1000ad, 'h1000d2, 'h1000ae, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h10003c, 'h2004f7, 'h1000dc, 'h1000dd, 'h1000de, 'h100047, 'h1000df, 'h1000af, 'h1000ab, 'h1000e0, 'h1000ac, 'h1000e1, 'h1000ad, 'h1000e2, 'h1000ae, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h10003c, 'h2004f7, 'h1000e9, 'h1000ea, 'h1000eb, 'h100047, 'h1000ec, 'h1000af, 'h1000ab, 'h1000ed, 'h1000ac, 'h1000ee, 'h1000ad, 'h1000ef, 'h1000ae, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h10003c, 'h2004f7, 'h1000f6, 'h1000f7, 'h1000f8, 'h100047, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000af, 'h1000fc, 'h1000ab, 'h1000ac, 'h1000fd, 'h1000ad, 'h1000fe, 'h1000ae, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h10003c, 'h2004f7, 'h100103, 'h100104, 'h100105, 'h100047, 'h100106, 'h100107, 'h100108, 'h1000af, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h1000ab, 'h1000ac, 'h10010d, 'h1000ad, 'h10010e, 'h1000ae, 'h10010f, 'h10003c, 'h2004f7, 'h100110, 'h100111, 'h100112, 'h100047, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h1000af, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h1000ab, 'h1000ac, 'h10011d, 'h1000ad, 'h10003c, 'h2004f7, 'h10011e, 'h1000ae, 'h10011f, 'h100047, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h1000af, 'h100125, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h1000ab, 'h10003c, 'h2004f7, 'h10012d, 'h1000ac, 'h10012e, 'h1000ad, 'h100047, 'h10012f, 'h1000ae, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h1000af, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h1000ab, 'h10003c, 'h2004f7, 'h10013a, 'h1000ac, 'h10013b, 'h1000ad, 'h100047, 'h10013c, 'h1000ae, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h1000af, 'h100145, 'h100146, 'h100147, 'h10003c, 'h2004f7, 'h100148, 'h1000ab, 'h100149, 'h1000ac, 'h100047, 'h10014a, 'h1000ad, 'h10014b, 'h1000ae, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h1000af, 'h10003c, 'h2004f7, 'h100155, 'h1000ab, 'h100156, 'h1000ac, 'h100047, 'h100157, 'h1000ad, 'h100158, 'h1000ae, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h10003c, 'h2004f7, 'h100163, 'h100164, 'h1000af, 'h1000ab, 'h100047, 'h100165, 'h1000ac, 'h100166, 'h1000ad, 'h100167, 'h1000ae, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h10003c, 'h2004f7, 'h100170, 'h1000b3, 'h1000af, 'h1000b4, 'h100047, 'h1000b0, 'h1000b5, 'h1000b1, 'h1000b6, 'h1000b2, 'h1000b7, 'h1000b8, 'h1000b9, 'h1000ba, 'h1000bb, 'h1000bc, 'h1000bd, 'h1000be, 'h1000bf, 'h10003c, 'h2004f7, 'h1000c0, 'h1000c1, 'h1000c2, 'h1000c3, 'h100047, 'h1000b3, 'h1000af, 'h1000c4, 'h1000b0, 'h1000c5, 'h1000b1, 'h1000c6, 'h1000b2, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h1000cc, 'h10003c, 'h2004f7, 'h1000cd, 'h1000ce, 'h1000cf, 'h1000d0, 'h100047, 'h1000d1, 'h1000d2, 'h1000d3, 'h1000b3, 'h1000af, 'h1000d4, 'h1000b0, 'h1000d5, 'h1000b1, 'h1000d6, 'h1000b2, 'h1000d7, 'h1000d8, 'h1000d9, 'h10003c, 'h2004f7, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h100047, 'h1000de, 'h1000df, 'h1000e0, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000b3, 'h1000e4, 'h1000af, 'h1000b0, 'h1000e5, 'h1000b1, 'h1000e6, 'h1000b2, 'h10003c, 'h2004f7, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h100047, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h1000f0, 'h1000b3, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000af, 'h1000b0, 'h1000f5, 'h10003c, 'h2004f7, 'h1000b1, 'h1000f6, 'h1000b2, 'h1000f7, 'h100047, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h1000b3, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h10003c, 'h2004f7, 'h1000af, 'h1000b0, 'h100105, 'h1000b1, 'h100047, 'h100106, 'h1000b2, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h1000b3, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h10003c, 'h2004f7, 'h100112, 'h100113, 'h100114, 'h1000af, 'h100047, 'h1000b0, 'h100115, 'h1000b1, 'h100116, 'h1000b2, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h1000b3, 'h10011c, 'h10011d, 'h10011e, 'h10003c, 'h2004f7, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100047, 'h100123, 'h100124, 'h1000af, 'h1000b0, 'h100125, 'h1000b1, 'h100126, 'h1000b2, 'h100127, 'h100128, 'h1000b3, 'h100129, 'h10012a, 'h10012b, 'h10003c, 'h2004f7, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100047, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h1000af, 'h100135, 'h1000b0, 'h100136, 'h1000b1, 'h100137, 'h1000b2, 'h100138, 'h1000b3, 'h10003c, 'h2004f7, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h100047, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h1000af, 'h100142, 'h1000b0, 'h100143, 'h1000b1, 'h100144, 'h1000b2, 'h100145, 'h100146, 'h10003c, 'h2004f7, 'h100147, 'h100148, 'h1000b3, 'h100149, 'h100047, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h1000af, 'h100151, 'h1000b0, 'h100152, 'h1000b1, 'h100153, 'h1000b2, 'h10003c, 'h2004f7, 'h100154, 'h100155, 'h100156, 'h100157, 'h100047, 'h100158, 'h1000b3, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h1000af, 'h10015e, 'h1000b0, 'h10015f, 'h1000b1, 'h100160, 'h1000b2, 'h10003c, 'h2004f7, 'h100161, 'h100162, 'h100163, 'h100164, 'h100047, 'h100165, 'h100166, 'h100167, 'h100168, 'h1000b3, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h1000af, 'h1000b0, 'h10016e, 'h1000b1, 'h10003c, 'h2004f7, 'h10016f, 'h1000b2, 'h100170, 'h1000b7, 'h1000ba, 'h100047, 'h1000b8, 'h1000b4, 'h1000b9, 'h1000b5, 'h1000b6, 'h1000bb, 'h1000be, 'h1000b3, 'h1000bc, 'h1000bd, 'h1000bf, 'h1000c3, 'h1000c0, 'h10003c, 'h2004f7, 'h1000c1, 'h1000c2, 'h1000c7, 'h1000b7, 'h1000c4, 'h100047, 'h1000c5, 'h1000b4, 'h1000c6, 'h1000b5, 'h1000b6, 'h1000cb, 'h1000c8, 'h1000b3, 'h1000c9, 'h1000ca, 'h1000cf, 'h1000cc, 'h1000cd, 'h10003c, 'h2004f7, 'h1000ce, 'h1000d3, 'h1000d0, 'h1000d1, 'h1000d2, 'h100047, 'h1000b7, 'h1000d7, 'h1000d4, 'h1000b4, 'h1000d5, 'h1000b5, 'h1000d6, 'h1000b6, 'h1000db, 'h1000b3, 'h1000d8, 'h1000d9, 'h1000da, 'h10003c, 'h2004f7, 'h1000df, 'h1000dc, 'h1000dd, 'h1000de, 'h1000e3, 'h100047, 'h1000b7, 'h1000e0, 'h1000e1, 'h1000b4, 'h1000e2, 'h1000b5, 'h1000e4, 'h1000e7, 'h1000e5, 'h1000e6, 'h1000b6, 'h1000e8, 'h1000eb, 'h10003c, 'h2004f7, 'h1000b3, 'h1000e9, 'h1000ea, 'h1000ec, 'h1000ef, 'h100047, 'h1000b7, 'h1000ed, 'h1000ee, 'h1000f0, 'h1000f3, 'h1000b4, 'h1000f1, 'h1000b5, 'h1000f2, 'h1000f4, 'h1000f7, 'h1000f5, 'h1000f6, 'h10003c, 'h2004f7, 'h1000b6, 'h1000f8, 'h1000fb, 'h1000b3, 'h1000f9, 'h100047, 'h1000fa, 'h1000b7, 'h1000fc, 'h1000ff, 'h1000fd, 'h1000b4, 'h1000fe, 'h1000b5, 'h100100, 'h100103, 'h100101, 'h100102, 'h100104, 'h100107, 'h10003c, 'h2004f7, 'h100105, 'h100106, 'h1000b6, 'h100108, 'h10010b, 'h100047, 'h1000b7, 'h1000b3, 'h100109, 'h10010a, 'h10010c, 'h10010f, 'h1000b4, 'h10010d, 'h1000b5, 'h10010e, 'h100110, 'h100113, 'h100111, 'h10003c, 'h2004f7, 'h100112, 'h100114, 'h100117, 'h100115, 'h100116, 'h100047, 'h1000b6, 'h1000b7, 'h100118, 'h10011b, 'h1000b3, 'h100119, 'h1000b4, 'h10011a, 'h1000b5, 'h10011c, 'h10011f, 'h10011d, 'h10011e, 'h10003c, 'h2004f7, 'h100120, 'h100123, 'h100121, 'h100122, 'h100124, 'h100127, 'h100047, 'h1000b7, 'h100125, 'h100126, 'h1000b6, 'h100128, 'h10012b, 'h1000b3, 'h1000b4, 'h100129, 'h1000b5, 'h10012a, 'h10012c, 'h10012f, 'h10003c, 'h2004f7, 'h10012d, 'h10012e, 'h100130, 'h100133, 'h100131, 'h100047, 'h100132, 'h1000b7, 'h100134, 'h100137, 'h100135, 'h100136, 'h1000b6, 'h100138, 'h10013b, 'h1000b3, 'h100139, 'h1000b4, 'h10013a, 'h10003c, 'h2004f7, 'h1000b5, 'h10013c, 'h10013f, 'h10013d, 'h10013e, 'h100047, 'h100140, 'h1000b7, 'h100144, 'h100141, 'h100142, 'h100143, 'h1000b6, 'h100148, 'h100145, 'h1000b3, 'h100146, 'h1000b4, 'h100147, 'h10003c, 'h2004f7, 'h1000b5, 'h10014c, 'h100149, 'h10014a, 'h10014b, 'h100047, 'h100150, 'h1000b7, 'h10014d, 'h10014e, 'h10014f, 'h100154, 'h100151, 'h100152, 'h100153, 'h1000b6, 'h100158, 'h1000b3, 'h100155, 'h10003c, 'h2004f7, 'h1000b4, 'h100156, 'h1000b5, 'h100157, 'h10015c, 'h100047, 'h100159, 'h10015a, 'h10015b, 'h1000b7, 'h100160, 'h10015d, 'h10015e, 'h10015f, 'h100164, 'h100161, 'h100162, 'h100163, 'h1000b6, 'h10003c, 'h2004f7, 'h100165, 'h100168, 'h1000b3, 'h1000b4, 'h100166, 'h100047, 'h1000b5, 'h100167, 'h100169, 'h1000b7, 'h10016c, 'h10016a, 'h10016b, 'h10016d, 'h100170, 'h10016e, 'h10016f, 'h1000bb, 'h1000bf, 'h10003c, 'h2004f7, 'h1000bc, 'h1000b8, 'h1000bd, 'h1000b9, 'h1000be, 'h100047, 'h1000ba, 'h1000c3, 'h1000c0, 'h1000b7, 'h1000c1, 'h1000c2, 'h1000c7, 'h1000c4, 'h1000c5, 'h1000c6, 'h1000cb, 'h1000bb, 'h1000c8, 'h10003c, 'h2004f7, 'h1000c9, 'h1000b8, 'h1000ca, 'h1000b9, 'h1000cf, 'h100047, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000ba, 'h1000d3, 'h1000b7, 'h1000d0, 'h1000d1, 'h1000d2, 'h1000d7, 'h1000d4, 'h1000d5, 'h1000d6, 'h10003c, 'h2004f7, 'h1000bb, 'h1000db, 'h1000d8, 'h1000b8, 'h1000d9, 'h100047, 'h1000b9, 'h1000da, 'h1000df, 'h1000dc, 'h1000dd, 'h1000de, 'h1000ba, 'h1000e0, 'h1000e3, 'h1000b7, 'h1000e1, 'h1000e2, 'h1000e4, 'h1000e7, 'h10003c, 'h2004f7, 'h1000bb, 'h1000e5, 'h1000b8, 'h1000e6, 'h100047, 'h1000b9, 'h1000e8, 'h1000eb, 'h1000e9, 'h1000ea, 'h1000ec, 'h1000ef, 'h1000ed, 'h1000ee, 'h1000ba, 'h1000f0, 'h1000f3, 'h1000b7, 'h1000f1, 'h10003c, 'h2004f7, 'h1000f2, 'h1000bb, 'h1000f4, 'h1000f7, 'h100047, 'h1000b8, 'h1000f5, 'h1000b9, 'h1000f6, 'h1000f8, 'h1000fb, 'h1000f9, 'h1000fa, 'h1000fc, 'h1000ff, 'h1000fd, 'h1000fe, 'h1000ba, 'h100100, 'h100103, 'h10003c, 'h2004f7, 'h1000bb, 'h1000b7, 'h100101, 'h100047, 'h1000b8, 'h100102, 'h1000b9, 'h100104, 'h100107, 'h100105, 'h100106, 'h100108, 'h10010b, 'h100109, 'h10010a, 'h10010c, 'h10010f, 'h10010d, 'h10010e, 'h10003c, 'h2004f7, 'h1000ba, 'h1000bb, 'h100110, 'h100113, 'h100047, 'h1000b7, 'h1000b8, 'h100111, 'h1000b9, 'h100112, 'h100114, 'h100117, 'h100115, 'h100116, 'h100118, 'h10011b, 'h100119, 'h10011a, 'h10011c, 'h10011f, 'h10003c, 'h2004f7, 'h1000bb, 'h10011d, 'h10011e, 'h100047, 'h1000ba, 'h100120, 'h100123, 'h1000b7, 'h1000b8, 'h100121, 'h1000b9, 'h100122, 'h100124, 'h100127, 'h100125, 'h100126, 'h100128, 'h10012b, 'h100129, 'h10003c, 'h2004f7, 'h10012a, 'h1000bb, 'h10012c, 'h10012f, 'h100047, 'h10012d, 'h10012e, 'h1000ba, 'h100130, 'h100133, 'h1000b7, 'h1000b8, 'h100131, 'h1000b9, 'h100132, 'h100134, 'h100137, 'h100135, 'h100136, 'h10003c, 'h2004f7, 'h100138, 'h1000bb, 'h10013b, 'h100139, 'h100047, 'h10013a, 'h10013c, 'h100140, 'h10013d, 'h10013e, 'h10013f, 'h1000ba, 'h100144, 'h1000b7, 'h100141, 'h1000b8, 'h100142, 'h1000b9, 'h100143, 'h10003c, 'h2004f7, 'h100148, 'h1000bb, 'h100145, 'h100146, 'h100047, 'h100147, 'h10014c, 'h100149, 'h10014a, 'h10014b, 'h100150, 'h10014d, 'h10014e, 'h10014f, 'h1000ba, 'h100154, 'h1000b7, 'h100151, 'h1000b8, 'h10003c, 'h2004f7, 'h100152, 'h1000b9, 'h100153, 'h1000bb, 'h100047, 'h100158, 'h100155, 'h100156, 'h100157, 'h10015c, 'h100159, 'h10015a, 'h10015b, 'h100160, 'h10015d, 'h10015e, 'h10015f, 'h1000ba, 'h100161, 'h100164, 'h10003c, 'h2004f7, 'h1000b7, 'h1000b8, 'h100162, 'h100047, 'h1000b9, 'h100163, 'h1000bb, 'h100165, 'h100168, 'h100166, 'h100167, 'h100169, 'h10016c, 'h10016a, 'h10016b, 'h10016d, 'h100170, 'h10016e, 'h10016f, 'h10003c, 'h2004f7, 'h1000ba, 'h1000bf, 'h1000c0, 'h100047, 'h1000bc, 'h1000c1, 'h1000bd, 'h1000c2, 'h1000be, 'h1000c3, 'h1000bb, 'h1000c4, 'h1000c5, 'h1000c6, 'h1000c7, 'h1000c8, 'h1000c9, 'h1000ca, 'h1000cb, 'h10003c, 'h2004f7, 'h1000cc, 'h1000cd, 'h1000ce, 'h100047, 'h1000cf, 'h1000bf, 'h1000d0, 'h1000bc, 'h1000d1, 'h1000bd, 'h1000d2, 'h1000be, 'h1000d3, 'h1000bb, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h10003c, 'h2004f7, 'h1000d9, 'h1000da, 'h1000db, 'h100047, 'h1000dc, 'h1000bf, 'h1000dd, 'h1000bc, 'h1000de, 'h1000bd, 'h1000df, 'h1000be, 'h1000e0, 'h1000bb, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h10003c, 'h2004f7, 'h1000e6, 'h1000e7, 'h1000e8, 'h100047, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000bf, 'h1000ec, 'h1000bc, 'h1000ed, 'h1000bd, 'h1000ee, 'h1000be, 'h1000ef, 'h1000f0, 'h1000bb, 'h1000f1, 'h1000f2, 'h10003c, 'h2004f7, 'h1000f3, 'h1000f4, 'h1000f5, 'h100047, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000bf, 'h1000f9, 'h1000bc, 'h1000fa, 'h1000bd, 'h1000fb, 'h1000be, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h10003c, 'h2004f7, 'h1000bb, 'h100101, 'h100102, 'h100047, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h1000bf, 'h100108, 'h1000bc, 'h100109, 'h1000bd, 'h10010a, 'h1000be, 'h10010b, 'h10010c, 'h10010d, 'h10003c, 'h2004f7, 'h10010e, 'h10010f, 'h100110, 'h100047, 'h1000bb, 'h100111, 'h100112, 'h100113, 'h100114, 'h1000bf, 'h100115, 'h1000bc, 'h100116, 'h1000bd, 'h100117, 'h1000be, 'h100118, 'h100119, 'h10011a, 'h10003c, 'h2004f7, 'h10011b, 'h10011c, 'h10011d, 'h100047, 'h10011e, 'h10011f, 'h100120, 'h1000bb, 'h100121, 'h100122, 'h100123, 'h1000bf, 'h100124, 'h1000bc, 'h100125, 'h1000bd, 'h100126, 'h1000be, 'h100127, 'h10003c, 'h2004f7, 'h100128, 'h100129, 'h10012a, 'h100047, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h1000bb, 'h100131, 'h100132, 'h100133, 'h1000bf, 'h100134, 'h1000bc, 'h100135, 'h1000bd, 'h10003c, 'h2004f7, 'h100136, 'h1000be, 'h100137, 'h100047, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h1000bb, 'h100141, 'h100142, 'h1000bc, 'h100143, 'h1000bd, 'h10003c, 'h2004f7, 'h100144, 'h1000be, 'h1000bf, 'h100047, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h1000bb, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h1000bc, 'h10003c, 'h2004f7, 'h100152, 'h1000bd, 'h100153, 'h100047, 'h1000be, 'h100154, 'h1000bf, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h1000bb, 'h10015e, 'h1000bc, 'h10003c, 'h2004f7, 'h10015f, 'h1000bd, 'h100160, 'h100047, 'h1000be, 'h100161, 'h1000bf, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10003c, 'h2004f7, 'h1000bb, 'h1000bc, 'h10016e, 'h100047, 'h1000bd, 'h10016f, 'h1000be, 'h100170, 'h1000bf, 'h1000c3, 'h1000c6, 'h1000c4, 'h1000c0, 'h1000c5, 'h1000c1, 'h1000c2, 'h1000c7, 'h1000ca, 'h1000c8, 'h10003c, 'h2004f7, 'h1000c9, 'h1000cb, 'h1000ce, 'h100047, 'h1000cc, 'h1000cd, 'h1000cf, 'h1000d2, 'h1000bf, 'h1000d0, 'h1000d1, 'h1000d3, 'h1000c3, 'h1000d6, 'h1000d4, 'h1000c0, 'h1000d5, 'h1000c1, 'h1000c2, 'h10003c, 'h2004f7, 'h1000d7, 'h1000d8, 'h1000da, 'h100047, 'h1000d9, 'h1000db, 'h1000dc, 'h1000de, 'h1000bf, 'h1000dd, 'h1000df, 'h1000e0, 'h1000c3, 'h1000e2, 'h1000e1, 'h1000c0, 'h1000e3, 'h1000e4, 'h1000e6, 'h10003c, 'h2004f7, 'h1000e5, 'h1000c1, 'h1000c2, 'h100047, 'h1000e7, 'h1000e8, 'h1000ea, 'h1000e9, 'h1000eb, 'h1000ec, 'h1000ee, 'h1000bf, 'h1000ed, 'h1000ef, 'h1000c3, 'h1000f0, 'h1000f2, 'h1000c0, 'h1000f1, 'h10003c, 'h2004f7, 'h1000f3, 'h1000f4, 'h1000f6, 'h100047, 'h1000f5, 'h1000c1, 'h1000c2, 'h1000f7, 'h1000f8, 'h1000fa, 'h1000f9, 'h1000fb, 'h1000fc, 'h1000fe, 'h1000c3, 'h1000bf, 'h1000fd, 'h1000c0, 'h1000ff, 'h10003c, 'h2004f7, 'h100100, 'h100102, 'h100101, 'h100047, 'h100103, 'h100104, 'h100106, 'h100105, 'h1000c1, 'h1000c2, 'h100107, 'h100108, 'h10010a, 'h100109, 'h10010b, 'h1000c3, 'h10010c, 'h10010e, 'h1000bf, 'h10003c, 'h2004f7, 'h1000c0, 'h10010d, 'h10010f, 'h100047, 'h100110, 'h100112, 'h100111, 'h100113, 'h100114, 'h100116, 'h100115, 'h1000c1, 'h1000c2, 'h100117, 'h100118, 'h1000c3, 'h10011b, 'h100119, 'h10011a, 'h10003c, 'h2004f7, 'h10011c, 'h10011f, 'h1000bf, 'h100047, 'h1000c0, 'h10011d, 'h10011e, 'h100120, 'h100123, 'h100121, 'h100122, 'h1000c1, 'h1000c2, 'h100124, 'h100127, 'h1000c3, 'h100125, 'h100126, 'h100128, 'h10012b, 'h10003c, 'h2004f7, 'h100129, 'h10012a, 'h100047, 'h10012c, 'h10012f, 'h1000bf, 'h1000c0, 'h10012d, 'h10012e, 'h100130, 'h100133, 'h100131, 'h1000c1, 'h100132, 'h1000c2, 'h1000c3, 'h100134, 'h100137, 'h100135, 'h10003c, 'h2004f7, 'h100136, 'h100138, 'h100047, 'h10013b, 'h100139, 'h10013a, 'h10013c, 'h10013f, 'h1000bf, 'h1000c0, 'h10013d, 'h10013e, 'h1000c1, 'h100140, 'h100143, 'h1000c3, 'h100141, 'h100142, 'h1000c2, 'h10003c, 'h2004f7, 'h100144, 'h100147, 'h100047, 'h100145, 'h100146, 'h100148, 'h10014b, 'h100149, 'h1000bf, 'h1000c0, 'h10014a, 'h10014c, 'h10014f, 'h10014d, 'h10014e, 'h1000c1, 'h100150, 'h1000c3, 'h100153, 'h10003c, 'h2004f7, 'h100151, 'h100152, 'h100047, 'h1000c2, 'h100154, 'h100157, 'h100155, 'h100156, 'h100158, 'h100159, 'h10015b, 'h1000bf, 'h1000c0, 'h10015a, 'h10015c, 'h10015d, 'h10015f, 'h1000c3, 'h10015e, 'h10003c, 'h2004f7, 'h1000c1, 'h100160, 'h100047, 'h1000c2, 'h100161, 'h100163, 'h100162, 'h100164, 'h100165, 'h100167, 'h100166, 'h100168, 'h100169, 'h10016b, 'h1000bf, 'h1000c0, 'h10016a, 'h10016c, 'h1000c3, 'h10003c, 'h2004f7, 'h10016d, 'h10016f, 'h100047, 'h10016e, 'h1000c1, 'h1000c2, 'h100170, 'h1000c7, 'h1000c8, 'h1000c4, 'h1000c9, 'h1000c5, 'h1000ca, 'h1000c6, 'h1000cb, 'h1000cc, 'h1000cd, 'h1000ce, 'h1000cf, 'h10003c, 'h2004f7, 'h1000d0, 'h1000c3, 'h100047, 'h1000d1, 'h1000d2, 'h1000d3, 'h1000d4, 'h1000c7, 'h1000d5, 'h1000c4, 'h1000d6, 'h1000c5, 'h1000d7, 'h1000c6, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h10003c, 'h2004f7, 'h1000dd, 'h1000de, 'h100047, 'h1000df, 'h1000e0, 'h1000c3, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000c7, 'h1000e4, 'h1000c4, 'h1000e5, 'h1000c5, 'h1000e6, 'h1000c6, 'h1000e7, 'h1000e8, 'h1000e9, 'h10003c, 'h2004f7, 'h1000ea, 'h1000eb, 'h100047, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h1000f0, 'h1000c3, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000c7, 'h1000f4, 'h1000c4, 'h1000f5, 'h1000c5, 'h1000f6, 'h1000c6, 'h10003c, 'h2004f7, 'h1000f7, 'h1000f8, 'h100047, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h1000c3, 'h100101, 'h100102, 'h100103, 'h1000c7, 'h100104, 'h1000c4, 'h100105, 'h10003c, 'h2004f7, 'h1000c5, 'h100106, 'h100047, 'h1000c6, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h1000c3, 'h100111, 'h100112, 'h100113, 'h1000c7, 'h10003c, 'h2004f7, 'h100114, 'h1000c4, 'h100047, 'h100115, 'h1000c5, 'h100116, 'h1000c6, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h1000c3, 'h100121, 'h10003c, 'h2004f7, 'h100122, 'h100123, 'h100047, 'h1000c7, 'h100124, 'h1000c4, 'h100125, 'h1000c5, 'h100126, 'h1000c6, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h10003c, 'h2004f7, 'h100130, 'h1000c3, 'h100047, 'h100131, 'h100132, 'h100133, 'h1000c7, 'h100134, 'h1000c4, 'h100135, 'h1000c5, 'h100136, 'h1000c6, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10003c, 'h2004f7, 'h10013d, 'h10013e, 'h100047, 'h10013f, 'h100140, 'h1000c3, 'h100141, 'h100142, 'h100143, 'h1000c7, 'h100144, 'h100145, 'h1000c4, 'h100146, 'h1000c5, 'h100147, 'h1000c6, 'h100148, 'h100149, 'h10003c, 'h2004f7, 'h10014a, 'h10014b, 'h100047, 'h10014c, 'h10014d, 'h1000c3, 'h10014e, 'h10014f, 'h100150, 'h1000c7, 'h100151, 'h100152, 'h1000c4, 'h100153, 'h1000c5, 'h100154, 'h1000c6, 'h100155, 'h100156, 'h10003c, 'h2004f7, 'h100157, 'h100158, 'h100047, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h1000c3, 'h10015e, 'h10015f, 'h100160, 'h1000c7, 'h100161, 'h1000c4, 'h100162, 'h1000c5, 'h100163, 'h1000c6, 'h10003c, 'h2004f7, 'h100164, 'h100165, 'h100047, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h1000c3, 'h10016e, 'h10016f, 'h100170, 'h1000c7, 'h1000cb, 'h1000cc, 'h1000c8, 'h10003c, 'h2004f7, 'h1000cd, 'h1000c9, 'h100047, 'h1000ce, 'h1000ca, 'h1000cf, 'h1000d0, 'h1000d1, 'h1000d2, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000c7, 'h1000d9, 'h1000da, 'h1000db, 'h10003c, 'h2004f7, 'h1000cb, 'h1000dc, 'h100047, 'h1000c8, 'h1000dd, 'h1000c9, 'h1000de, 'h1000ca, 'h1000df, 'h1000e0, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000c7, 'h10003c, 'h2004f7, 'h1000e9, 'h1000ea, 'h100047, 'h1000eb, 'h1000cb, 'h1000ec, 'h1000c8, 'h1000ed, 'h1000c9, 'h1000ee, 'h1000ca, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h10003c, 'h2004f7, 'h1000f7, 'h1000f8, 'h100047, 'h1000c7, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000cb, 'h1000fc, 'h1000c8, 'h1000fd, 'h1000c9, 'h1000fe, 'h1000ca, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h10003c, 'h2004f7, 'h100104, 'h100105, 'h100047, 'h100106, 'h100107, 'h100108, 'h1000c7, 'h100109, 'h10010a, 'h10010b, 'h1000cb, 'h10010c, 'h1000c8, 'h10010d, 'h1000c9, 'h10010e, 'h1000ca, 'h10010f, 'h100110, 'h10003c, 'h2004f7, 'h100111, 'h100112, 'h100047, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h1000c7, 'h100119, 'h10011a, 'h10011b, 'h1000cb, 'h10011c, 'h1000c8, 'h10011d, 'h1000c9, 'h10011e, 'h10003c, 'h2004f7, 'h1000ca, 'h10011f, 'h100047, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h1000c7, 'h100129, 'h10012a, 'h10012b, 'h1000cb, 'h10012c, 'h1000c8, 'h10003c, 'h2004f7, 'h10012d, 'h1000c9, 'h100047, 'h10012e, 'h1000ca, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h1000c7, 'h100139, 'h10013a, 'h10013b, 'h10003c, 'h2004f7, 'h1000cb, 'h10013c, 'h100047, 'h1000c8, 'h10013d, 'h1000c9, 'h10013e, 'h1000ca, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h1000c7, 'h10003c, 'h2004f7, 'h100149, 'h10014a, 'h100047, 'h10014b, 'h10014c, 'h1000cb, 'h10014d, 'h1000c8, 'h10014e, 'h1000c9, 'h10014f, 'h1000ca, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h1000c7, 'h10003c, 'h2004f7, 'h100156, 'h100157, 'h100047, 'h100158, 'h100159, 'h1000cb, 'h10015a, 'h1000c8, 'h10015b, 'h1000c9, 'h10015c, 'h1000ca, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h10003c, 'h2004f7, 'h100164, 'h100165, 'h100047, 'h1000c7, 'h100166, 'h100167, 'h100168, 'h1000cb, 'h100169, 'h1000c8, 'h10016a, 'h1000c9, 'h10016b, 'h1000ca, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h10003c, 'h2004f7, 'h1000d0, 'h1000cf, 'h100047, 'h1000cc, 'h1000d1, 'h1000cd, 'h1000d2, 'h1000ce, 'h1000d3, 'h1000d4, 'h1000d5, 'h1000d6, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h10003c, 'h2004f7, 'h1000de, 'h1000df, 'h100047, 'h1000cf, 'h1000e0, 'h1000cc, 'h1000e1, 'h1000cd, 'h1000e2, 'h1000ce, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h10003c, 'h2004f7, 'h1000ec, 'h1000ed, 'h100047, 'h1000ee, 'h1000ef, 'h1000cf, 'h1000f0, 'h1000cc, 'h1000f1, 'h1000cd, 'h1000f2, 'h1000ce, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h10003c, 'h2004f7, 'h1000fa, 'h1000fb, 'h100047, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h1000cf, 'h100100, 'h1000cc, 'h100101, 'h1000cd, 'h100102, 'h1000ce, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h10003c, 'h2004f7, 'h100108, 'h100109, 'h100047, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h1000cf, 'h100110, 'h1000cc, 'h100111, 'h1000cd, 'h100112, 'h1000ce, 'h100113, 'h100114, 'h100115, 'h10003c, 'h2004f7, 'h100116, 'h100117, 'h100047, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h1000cf, 'h100120, 'h1000cc, 'h100121, 'h1000cd, 'h100122, 'h1000ce, 'h100123, 'h10003c, 'h2004f7, 'h100124, 'h100125, 'h100047, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h1000cf, 'h100130, 'h1000cc, 'h100131, 'h1000cd, 'h100132, 'h10003c, 'h2004f7, 'h1000ce, 'h100133, 'h100047, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h1000cf, 'h100140, 'h1000cc, 'h100141, 'h10003c, 'h2004f7, 'h1000cd, 'h100142, 'h100047, 'h1000ce, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h1000cf, 'h10014e, 'h10014f, 'h100150, 'h10003c, 'h2004f7, 'h100151, 'h1000cc, 'h100047, 'h100152, 'h1000cd, 'h100153, 'h1000ce, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h1000cf, 'h10015d, 'h10015e, 'h10003c, 'h2004f7, 'h10015f, 'h100160, 'h100047, 'h100161, 'h1000cc, 'h100162, 'h1000cd, 'h100163, 'h1000ce, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h1000cf, 'h10003c, 'h2004f7, 'h10016d, 'h10016e, 'h100047, 'h10016f, 'h100170, 'h1000d4, 'h1000d3, 'h1000d0, 'h1000d5, 'h1000d1, 'h1000d6, 'h1000d2, 'h1000d7, 'h1000d8, 'h1000d9, 'h1000da, 'h1000db, 'h1000dc, 'h1000dd, 'h10003c, 'h2004f7, 'h1000de, 'h1000df, 'h100047, 'h1000e0, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000d3, 'h1000e4, 'h1000d0, 'h1000e5, 'h1000d1, 'h1000e6, 'h1000d2, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h10003c, 'h2004f7, 'h1000ec, 'h1000ed, 'h100047, 'h1000ee, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000d3, 'h1000f4, 'h1000d0, 'h1000f5, 'h1000d1, 'h1000f6, 'h1000d2, 'h1000f7, 'h1000f8, 'h1000f9, 'h10003c, 'h2004f7, 'h1000fa, 'h1000fb, 'h100047, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h1000d3, 'h100104, 'h1000d0, 'h100105, 'h1000d1, 'h100106, 'h1000d2, 'h100107, 'h10003c, 'h2004f7, 'h100108, 'h100109, 'h100047, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h1000d3, 'h100114, 'h1000d0, 'h100115, 'h1000d1, 'h100116, 'h10003c, 'h2004f7, 'h1000d2, 'h100117, 'h100047, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h1000d3, 'h100124, 'h1000d0, 'h100125, 'h10003c, 'h2004f7, 'h1000d1, 'h100126, 'h100047, 'h1000d2, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h1000d3, 'h100134, 'h10003c, 'h2004f7, 'h1000d0, 'h100135, 'h100047, 'h1000d1, 'h100136, 'h1000d2, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h10003c, 'h2004f7, 'h1000d3, 'h100144, 'h100047, 'h100145, 'h1000d0, 'h1000d1, 'h100146, 'h1000d2, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h10003c, 'h2004f7, 'h1000d3, 'h100152, 'h100047, 'h100153};
	
endpackage
