

package LU_PKG_3;
	
	import LU_PKG_2::DATA2;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h10026c, 'h2004f8, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100170, 'h10009e, 'h10003c, 'h100047, 'h10009b, 'h100171, 'h10009c, 'h100172, 'h10009d, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h2004f8, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h10009e, 'h100180, 'h100181, 'h10009b, 'h10009c, 'h100182, 'h10009d, 'h100183, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h10009e, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h10009b, 'h10009c, 'h100192, 'h10009d, 'h100193, 'h2004f8, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h10009e, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h10009b, 'h1001a2, 'h10009c, 'h2004f8, 'h1001a3, 'h10009d, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h10009e, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h10009b, 'h2004f8, 'h1001b2, 'h10009c, 'h1001b3, 'h10009d, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h100047, 'h1001b8, 'h10009e, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h2004f8, 'h1001c1, 'h10009b, 'h1001c2, 'h10009c, 'h1001c3, 'h10009d, 'h1001c4, 'h1001c5, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h10009e, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h2004f8, 'h1001cf, 'h1001d0, 'h1001d1, 'h10009b, 'h1001d2, 'h10009c, 'h1001d3, 'h10009d, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h10009e, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h2004f8, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h10009b, 'h1001e2, 'h10009c, 'h10003c, 'h100047, 'h1001e3, 'h10009d, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h10009e, 'h1001e9, 'h1001ea, 'h2004f8, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h10009b, 'h10003c, 'h100047, 'h1001f2, 'h10009c, 'h1001f3, 'h10009d, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h10009e, 'h2004f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h10003c, 'h100047, 'h100201, 'h100202, 'h10009b, 'h10009c, 'h100203, 'h10009d, 'h100204, 'h100205, 'h100206, 'h10009e, 'h2004f8, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10003c, 'h100047, 'h10020f, 'h100210, 'h100211, 'h100212, 'h10009b, 'h10009c, 'h100213, 'h10009d, 'h100214, 'h10009e, 'h2004f8, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10003c, 'h100047, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h10009b, 'h100223, 'h10009c, 'h100224, 'h2004f8, 'h10009d, 'h100225, 'h10009e, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10003c, 'h100047, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h10009b, 'h100233, 'h2004f8, 'h10009c, 'h100234, 'h10009d, 'h100235, 'h10009e, 'h100236, 'h100237, 'h100238, 'h10003c, 'h100047, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h2004f8, 'h10009b, 'h100243, 'h10009c, 'h100244, 'h10009d, 'h100245, 'h10009e, 'h100246, 'h10003c, 'h100047, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h2004f8, 'h100251, 'h100252, 'h10009b, 'h100253, 'h10009c, 'h100254, 'h10009d, 'h100255, 'h10003c, 'h100047, 'h10009e, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h2004f8, 'h10025f, 'h100260, 'h100261, 'h100262, 'h10009b, 'h100263, 'h10009c, 'h100264, 'h10003c, 'h100047, 'h10009d, 'h100265, 'h10009e, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h2004f8, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100170, 'h1000a2, 'h10003c, 'h100047, 'h10009f, 'h100171, 'h1000a0, 'h100172, 'h1000a1, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h2004f8, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h1000a2, 'h100180, 'h100181, 'h10009f, 'h1000a0, 'h100182, 'h1000a1, 'h100183, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h1000a2, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h10009f, 'h1000a0, 'h100192, 'h1000a1, 'h100193, 'h2004f8, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h1000a2, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h10009f, 'h1001a2, 'h1000a0, 'h2004f8, 'h1001a3, 'h1000a1, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h1000a2, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h10009f, 'h2004f8, 'h1001b2, 'h1000a0, 'h1001b3, 'h1000a1, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h100047, 'h1001b8, 'h1000a2, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h2004f8, 'h1001c1, 'h10009f, 'h1001c2, 'h1000a0, 'h1001c3, 'h1000a1, 'h1001c4, 'h1001c5, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1000a2, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h2004f8, 'h1001cf, 'h1001d0, 'h1001d1, 'h10009f, 'h1001d2, 'h1000a0, 'h1001d3, 'h1000a1, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1000a2, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h2004f8, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h10009f, 'h1001e2, 'h1000a0, 'h10003c, 'h100047, 'h1001e3, 'h1000a1, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1000a2, 'h1001e9, 'h1001ea, 'h2004f8, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h10009f, 'h10003c, 'h100047, 'h1001f2, 'h1000a0, 'h1001f3, 'h1000a1, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1000a2, 'h2004f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h10003c, 'h100047, 'h100201, 'h100202, 'h10009f, 'h1000a0, 'h100203, 'h1000a1, 'h100204, 'h100205, 'h100206, 'h1000a2, 'h2004f8, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10003c, 'h100047, 'h10020f, 'h100210, 'h100211, 'h100212, 'h10009f, 'h1000a0, 'h100213, 'h1000a1, 'h100214, 'h1000a2, 'h2004f8, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10003c, 'h100047, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h10009f, 'h100223, 'h1000a0, 'h100224, 'h1000a1, 'h2004f8, 'h100225, 'h1000a2, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10003c, 'h100047, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h10009f, 'h100233, 'h1000a0, 'h2004f8, 'h100234, 'h1000a1, 'h100235, 'h1000a2, 'h100236, 'h100237, 'h100238, 'h10003c, 'h100047, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h10009f, 'h2004f8, 'h100243, 'h1000a0, 'h100244, 'h1000a1, 'h100245, 'h1000a2, 'h100246, 'h10003c, 'h100047, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h2004f8, 'h100252, 'h10009f, 'h100253, 'h1000a0, 'h100254, 'h1000a1, 'h100255, 'h10003c, 'h100047, 'h1000a2, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h2004f8, 'h100260, 'h100261, 'h100262, 'h10009f, 'h100263, 'h1000a0, 'h100264, 'h10003c, 'h100047, 'h1000a1, 'h100265, 'h1000a2, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h2004f8, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100170, 'h1000a6, 'h10003c, 'h100047, 'h100171, 'h1000a3, 'h1000a4, 'h100172, 'h1000a5, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h2004f8, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h1000a6, 'h100180, 'h100181, 'h1000a3, 'h1000a4, 'h100182, 'h1000a5, 'h100183, 'h100184, 'h100185, 'h100186, 'h2004f8, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h1000a6, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h1000a3, 'h1000a4, 'h100192, 'h1000a5, 'h100193, 'h100194, 'h2004f8, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h1000a6, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h1000a3, 'h1000a4, 'h1001a2, 'h1000a5, 'h2004f8, 'h1001a3, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h1000a6, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1000a3, 'h1001b2, 'h2004f8, 'h1000a4, 'h1001b3, 'h1000a5, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h100047, 'h1001b8, 'h1000a6, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h2004f8, 'h1000a3, 'h1001c2, 'h1000a4, 'h1001c3, 'h1000a5, 'h1001c4, 'h1001c5, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1000a6, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h2004f8, 'h1001d0, 'h1001d1, 'h1000a3, 'h1001d2, 'h1000a4, 'h1001d3, 'h1000a5, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1000a6, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h2004f8, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1000a3, 'h1001e2, 'h1000a4, 'h10003c, 'h100047, 'h1001e3, 'h1000a5, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1000a6, 'h1001e9, 'h1001ea, 'h1001eb, 'h2004f8, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000a3, 'h10003c, 'h100047, 'h1000a4, 'h1001f3, 'h1000a5, 'h1001f4, 'h1001f5, 'h1001f6, 'h1000a6, 'h1001f7, 'h1001f8, 'h1001f9, 'h2004f8, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h10003c, 'h100047, 'h100202, 'h1000a3, 'h1000a4, 'h100203, 'h1000a5, 'h100204, 'h1000a6, 'h100205, 'h100206, 'h100207, 'h2004f8, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h10003c, 'h100047, 'h100210, 'h100211, 'h100212, 'h1000a3, 'h1000a4, 'h100213, 'h1000a5, 'h100214, 'h1000a6, 'h100215, 'h2004f8, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10003c, 'h100047, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000a3, 'h1000a4, 'h100223, 'h1000a5, 'h100224, 'h2004f8, 'h1000a6, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10003c, 'h100047, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h1000a3, 'h100233, 'h1000a4, 'h2004f8, 'h100234, 'h1000a5, 'h100235, 'h1000a6, 'h100236, 'h100237, 'h100238, 'h100239, 'h10003c, 'h100047, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h1000a3, 'h2004f8, 'h100243, 'h1000a4, 'h100244, 'h1000a5, 'h100245, 'h1000a6, 'h100246, 'h100247, 'h10003c, 'h100047, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h2004f8, 'h100252, 'h1000a3, 'h100253, 'h1000a4, 'h100254, 'h1000a5, 'h100255, 'h1000a6, 'h10003c, 'h100047, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h2004f8, 'h100260, 'h100261, 'h100262, 'h1000a3, 'h100263, 'h1000a4, 'h100264, 'h1000a5, 'h10003c, 'h100047, 'h100265, 'h1000a6, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h2004f8, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000ab, 'h1000a7, 'h10003c, 'h100047, 'h1000a8, 'h100172, 'h1000a9, 'h100173, 'h1000aa, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h2004f8, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h10003c, 'h100047, 'h100181, 'h1000ab, 'h1000a7, 'h1000a8, 'h100182, 'h1000a9, 'h100183, 'h1000aa, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h1000ab, 'h1000a7, 'h1000a8, 'h100192, 'h1000a9, 'h100193, 'h2004f8, 'h1000aa, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10003c, 'h100047, 'h10019b, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h1000ab, 'h1000a7, 'h1000a8, 'h2004f8, 'h1001a2, 'h1000a9, 'h1001a3, 'h1000aa, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h10003c, 'h100047, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h2004f8, 'h1000ab, 'h1000a7, 'h1001b2, 'h1000a8, 'h1001b3, 'h1000a9, 'h1001b4, 'h1000aa, 'h10003c, 'h100047, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h2004f8, 'h1001bf, 'h1001c0, 'h1001c1, 'h1000ab, 'h1000a7, 'h1001c2, 'h1000a8, 'h1001c3, 'h10003c, 'h100047, 'h1000a9, 'h1001c4, 'h1000aa, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h2004f8, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1000ab, 'h1000a7, 'h10003c, 'h100047, 'h1001d2, 'h1000a8, 'h1001d3, 'h1000a9, 'h1001d4, 'h1000aa, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h2004f8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1000ab, 'h1000a7, 'h10003c, 'h100047, 'h1001df, 'h1000a8, 'h1001e0, 'h1000a9, 'h1001e1, 'h1000aa, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h2004f8, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h10003c, 'h100047, 'h1000ab, 'h1001ee, 'h1000a7, 'h1000a8, 'h1001ef, 'h1000a9, 'h1001f0, 'h1000aa, 'h1001f1, 'h1001f2, 'h2004f8, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h10003c, 'h100047, 'h1000ab, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1000a7, 'h1000a8, 'h1001ff, 'h1000a9, 'h100200, 'h2004f8, 'h1000aa, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100207, 'h10003c, 'h100047, 'h100208, 'h100209, 'h10020a, 'h1000ab, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h1000a7, 'h1000a8, 'h2004f8, 'h10020f, 'h1000a9, 'h100210, 'h1000aa, 'h100211, 'h100212, 'h100213, 'h100214, 'h10003c, 'h100047, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h1000ab, 'h10021b, 'h10021c, 'h10021d, 'h2004f8, 'h10021e, 'h1000a7, 'h1000a8, 'h10021f, 'h1000a9, 'h100220, 'h1000aa, 'h100221, 'h10003c, 'h100047, 'h100222, 'h100223, 'h100224, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h1000ab, 'h2004f8, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h1000a7, 'h10022f, 'h1000a8, 'h100230, 'h10003c, 'h100047, 'h1000a9, 'h100231, 'h1000aa, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h2004f8, 'h100239, 'h10023a, 'h1000ab, 'h10023b, 'h1000a7, 'h10023c, 'h1000a8, 'h10023d, 'h10003c, 'h100047, 'h1000a9, 'h10023e, 'h1000aa, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h2004f8, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h1000ab, 'h1000a7, 'h10024b, 'h10003c, 'h100047, 'h1000a8, 'h10024c, 'h1000a9, 'h10024d, 'h1000aa, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h2004f8, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10003c, 'h100047, 'h1000ab, 'h10025b, 'h1000a7, 'h1000a8, 'h10025c, 'h1000a9, 'h10025d, 'h1000aa, 'h10025e, 'h10025f, 'h2004f8, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h10003c, 'h100047, 'h1000ab, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h1000a7, 'h1000a8, 'h10026c, 'h1000a9, 'h10026d, 'h2004f8, 'h1000aa, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000af, 'h10003c, 'h100047, 'h1000ab, 'h1000ac, 'h100172, 'h1000ad, 'h100173, 'h1000ae, 'h100174, 'h100175, 'h100176, 'h100177, 'h2004f8, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h100180, 'h1000af, 'h100181, 'h1000ab, 'h1000ac, 'h100182, 'h1000ad, 'h100183, 'h1000ae, 'h100184, 'h2004f8, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10003c, 'h100047, 'h10018d, 'h1000af, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h1000ab, 'h1000ac, 'h100192, 'h1000ad, 'h2004f8, 'h100193, 'h1000ae, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10003c, 'h100047, 'h10019a, 'h10019b, 'h10019c, 'h1000af, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h1000ab, 'h2004f8, 'h1000ac, 'h1001a2, 'h1000ad, 'h1001a3, 'h1000ae, 'h1001a4, 'h1001a5, 'h1001a6, 'h10003c, 'h100047, 'h1001a7, 'h1001a8, 'h1001a9, 'h1000af, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h2004f8, 'h1001b0, 'h1001b1, 'h1000ab, 'h1001b2, 'h1000ac, 'h1001b3, 'h1000ad, 'h1001b4, 'h10003c, 'h100047, 'h1000ae, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1000af, 'h1001ba, 'h1001bb, 'h1001bc, 'h2004f8, 'h1001bd, 'h1001be, 'h1000ab, 'h1001bf, 'h1000ac, 'h1001c0, 'h1000ad, 'h1001c1, 'h10003c, 'h100047, 'h1000ae, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1000af, 'h2004f8, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1000ab, 'h1001ce, 'h1000ac, 'h1001cf, 'h10003c, 'h100047, 'h1000ad, 'h1001d0, 'h1000ae, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h2004f8, 'h1001d8, 'h1001d9, 'h1000af, 'h1001da, 'h1000ab, 'h1001db, 'h1000ac, 'h1001dc, 'h10003c, 'h100047, 'h1000ad, 'h1001dd, 'h1000ae, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h2004f8, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1000af, 'h1001ea, 'h1000ab, 'h10003c, 'h100047, 'h1000ac, 'h1001eb, 'h1000ad, 'h1001ec, 'h1000ae, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h2004f8, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1000af, 'h1001f7, 'h1001f8, 'h10003c, 'h100047, 'h1001f9, 'h1001fa, 'h1000ab, 'h1000ac, 'h1001fb, 'h1000ad, 'h1001fc, 'h1000ae, 'h1001fd, 'h1001fe, 'h2004f8, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h1000af, 'h10003c, 'h100047, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h1000ab, 'h1000ac, 'h10020b, 'h1000ad, 'h10020c, 'h2004f8, 'h1000ae, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000af, 'h10003c, 'h100047, 'h100213, 'h100214, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h1000ab, 'h1000ac, 'h2004f8, 'h10021b, 'h1000ad, 'h10021c, 'h1000ae, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h10003c, 'h100047, 'h100221, 'h1000af, 'h100222, 'h100223, 'h100224, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h2004f8, 'h10022a, 'h1000ab, 'h1000ac, 'h10022b, 'h1000ad, 'h10022c, 'h1000ae, 'h10022d, 'h10003c, 'h100047, 'h10022e, 'h1000af, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h2004f8, 'h100237, 'h1000ab, 'h1000ac, 'h100238, 'h1000ad, 'h100239, 'h1000ae, 'h10023a, 'h10003c, 'h100047, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h1000af, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h2004f8, 'h100244, 'h100245, 'h100246, 'h1000ab, 'h100247, 'h1000ac, 'h100248, 'h1000ad, 'h10003c, 'h100047, 'h100249, 'h1000ae, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h1000af, 'h10024f, 'h100250, 'h2004f8, 'h100251, 'h100252, 'h100253, 'h1000ab, 'h100254, 'h1000ac, 'h100255, 'h1000ad, 'h10003c, 'h100047, 'h100256, 'h1000ae, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h2004f8, 'h1000af, 'h10025f, 'h100260, 'h100261, 'h100262, 'h1000ab, 'h100263, 'h1000ac, 'h10003c, 'h100047, 'h100264, 'h1000ad, 'h100265, 'h1000ae, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h2004f8, 'h10026c, 'h10026d, 'h10026e, 'h1000af, 'h10026f, 'h1000ab, 'h100270, 'h1000ac, 'h10003c, 'h100047, 'h100271, 'h1000ad, 'h100272, 'h1000ae, 'h100171, 'h1000b3, 'h1000b0, 'h100172, 'h1000b1, 'h100173, 'h2004f8, 'h1000b2, 'h100174, 'h100175, 'h1000af, 'h100176, 'h100177, 'h100178, 'h100179, 'h10003c, 'h100047, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000b3, 'h100181, 'h1000b0, 'h2004f8, 'h100182, 'h1000b1, 'h100183, 'h1000b2, 'h100184, 'h100185, 'h1000af, 'h100186, 'h10003c, 'h100047, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h1000b3, 'h10018e, 'h1000b0, 'h2004f8, 'h10018f, 'h1000b1, 'h100190, 'h1000b2, 'h100191, 'h100192, 'h100193, 'h100194, 'h10003c, 'h100047, 'h100195, 'h1000af, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h1000b3, 'h2004f8, 'h10019d, 'h1000b0, 'h10019e, 'h1000b1, 'h10019f, 'h1000b2, 'h1001a0, 'h1001a1, 'h10003c, 'h100047, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1000af, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1000b3, 'h2004f8, 'h1001aa, 'h1000b0, 'h1001ab, 'h1000b1, 'h1001ac, 'h1000b2, 'h1001ad, 'h1001ae, 'h10003c, 'h100047, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1000af, 'h1001b6, 'h1001b7, 'h2004f8, 'h1001b8, 'h1001b9, 'h1000b3, 'h1001ba, 'h1000b0, 'h1001bb, 'h1000b1, 'h1001bc, 'h10003c, 'h100047, 'h1000b2, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1000af, 'h1001c3, 'h1001c4, 'h2004f8, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1000b3, 'h1001ca, 'h1000b0, 'h10003c, 'h100047, 'h1001cb, 'h1000b1, 'h1001cc, 'h1000b2, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1000af, 'h2004f8, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h10003c, 'h100047, 'h1000b3, 'h1001da, 'h1000b0, 'h1001db, 'h1000b1, 'h1001dc, 'h1000b2, 'h1001dd, 'h1001de, 'h1000af, 'h2004f8, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h10003c, 'h100047, 'h1001e7, 'h1001e8, 'h1001e9, 'h1000b3, 'h1001ea, 'h1000b0, 'h1001eb, 'h1000b1, 'h1001ec, 'h1000b2, 'h2004f8, 'h1001ed, 'h1001ee, 'h1000af, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h10003c, 'h100047, 'h1001f4, 'h1001f5, 'h1001f6, 'h1000b3, 'h1001f7, 'h1000b0, 'h1001f8, 'h1000b1, 'h1001f9, 'h1000b2, 'h2004f8, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1000af, 'h1001ff, 'h100200, 'h10003c, 'h100047, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h1000b3, 'h100206, 'h1000b0, 'h100207, 'h1000b1, 'h2004f8, 'h100208, 'h1000b2, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10003c, 'h100047, 'h1000af, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000b3, 'h100213, 'h1000b0, 'h100214, 'h1000b1, 'h2004f8, 'h100215, 'h1000b2, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10003c, 'h100047, 'h10021c, 'h10021d, 'h10021e, 'h1000af, 'h10021f, 'h100220, 'h100221, 'h1000b3, 'h100222, 'h1000b0, 'h2004f8, 'h100223, 'h1000b1, 'h100224, 'h1000b2, 'h100225, 'h100226, 'h100227, 'h100228, 'h10003c, 'h100047, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h1000af, 'h10022f, 'h100230, 'h100231, 'h2004f8, 'h1000b3, 'h100232, 'h100233, 'h1000b0, 'h100234, 'h1000b1, 'h100235, 'h1000b2, 'h10003c, 'h100047, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h1000af, 'h10023c, 'h10023d, 'h10023e, 'h2004f8, 'h1000b3, 'h10023f, 'h100240, 'h1000b0, 'h100241, 'h1000b1, 'h100242, 'h1000b2, 'h10003c, 'h100047, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h1000af, 'h10024b, 'h2004f8, 'h10024c, 'h10024d, 'h10024e, 'h1000b3, 'h10024f, 'h1000b0, 'h100250, 'h1000b1, 'h10003c, 'h100047, 'h100251, 'h1000b2, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h1000af, 'h100258, 'h2004f8, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h1000b3, 'h10025f, 'h10003c, 'h100047, 'h1000b0, 'h100260, 'h1000b1, 'h100261, 'h1000b2, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h2004f8, 'h100267, 'h1000af, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h1000b3, 'h10026c, 'h10003c, 'h100047, 'h1000b0, 'h10026d, 'h1000b1, 'h10026e, 'h1000b2, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h2004f8, 'h1000b7, 'h100174, 'h1000b4, 'h100172, 'h1000b5, 'h100173, 'h1000b6, 'h100175, 'h100178, 'h10003c, 'h100047, 'h1000b3, 'h100176, 'h100177, 'h100179, 'h10017c, 'h10017a, 'h10017b, 'h10017d, 'h100180, 'h2004f8, 'h1000b7, 'h10017e, 'h1000b4, 'h10017f, 'h1000b5, 'h100181, 'h100184, 'h100182, 'h100183, 'h10003c, 'h100047, 'h1000b6, 'h100185, 'h100188, 'h1000b3, 'h100186, 'h100187, 'h100189, 'h10018c, 'h10018a, 'h2004f8, 'h10018b, 'h1000b7, 'h10018d, 'h100190, 'h1000b4, 'h10018e, 'h1000b5, 'h10018f, 'h100191, 'h100194, 'h10003c, 'h100047, 'h100192, 'h100193, 'h1000b6, 'h100195, 'h100198, 'h1000b3, 'h100196, 'h100197, 'h2004f8, 'h100199, 'h1000b7, 'h10019c, 'h10019a, 'h1000b4, 'h10019b, 'h1000b5, 'h10019d, 'h1001a0, 'h10019e, 'h10003c, 'h100047, 'h10019f, 'h1001a1, 'h1001a4, 'h1001a2, 'h1001a3, 'h1000b6, 'h1001a5, 'h1001a8, 'h2004f8, 'h1000b3, 'h1001a6, 'h1001a7, 'h1000b7, 'h1001a9, 'h1001ac, 'h1000b4, 'h1001aa, 'h1000b5, 'h1001ab, 'h10003c, 'h100047, 'h1001ad, 'h1001b0, 'h1001ae, 'h1001af, 'h1001b1, 'h1001b4, 'h1001b2, 'h1001b3, 'h2004f8, 'h1000b6, 'h1001b5, 'h1001b8, 'h1000b7, 'h1000b3, 'h1001b6, 'h1000b4, 'h1001b7, 'h1000b5, 'h1001b9, 'h10003c, 'h100047, 'h1001bc, 'h1001ba, 'h1001bb, 'h1001bd, 'h1001c0, 'h1001be, 'h1001bf, 'h1001c1, 'h2004f8, 'h1000b6, 'h1001c5, 'h1001c2, 'h1001c3, 'h1001c4, 'h1000b7, 'h1001c9, 'h1000b3, 'h1001c6, 'h1000b4, 'h10003c, 'h100047, 'h1001c7, 'h1000b5, 'h1001c8, 'h1001cd, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001d1, 'h2004f8, 'h1001ce, 'h1001cf, 'h1001d0, 'h1000b6, 'h1001d5, 'h1000b7, 'h1001d2, 'h1000b3, 'h1001d3, 'h1000b4, 'h10003c, 'h100047, 'h1001d4, 'h1000b5, 'h1001d9, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001dd, 'h1001da, 'h2004f8, 'h1001db, 'h1001dc, 'h1001e1, 'h1001de, 'h1001df, 'h1001e0, 'h1000b6, 'h1000b7, 'h1001e5, 'h1001e2, 'h1000b3, 'h10003c, 'h100047, 'h1000b4, 'h1001e3, 'h1000b5, 'h1001e4, 'h1001e6, 'h1001e9, 'h1001e7, 'h2004f8, 'h1001e8, 'h1001ea, 'h1001ed, 'h1001eb, 'h1001ec, 'h1001ee, 'h1001f1, 'h1000b7, 'h1001ef, 'h1001f0, 'h1000b6, 'h10003c, 'h100047, 'h1001f2, 'h1001f5, 'h1000b3, 'h1000b4, 'h1001f3, 'h1000b5, 'h1001f4, 'h2004f8, 'h1001f6, 'h1001f9, 'h1001f7, 'h1001f8, 'h1001fa, 'h1001fd, 'h1001fb, 'h1001fc, 'h1000b7, 'h1001fe, 'h100201, 'h10003c, 'h100047, 'h1001ff, 'h100200, 'h1000b6, 'h100202, 'h100205, 'h1000b3, 'h1000b4, 'h2004f8, 'h100203, 'h1000b5, 'h100204, 'h100206, 'h100209, 'h100207, 'h100208, 'h10020a, 'h1000b7, 'h10020d, 'h10020b, 'h10003c, 'h100047, 'h10020c, 'h10020e, 'h100211, 'h10020f, 'h100210, 'h1000b6, 'h100212, 'h2004f8, 'h100215, 'h1000b3, 'h1000b4, 'h100213, 'h1000b5, 'h100214, 'h100216, 'h100219, 'h1000b7, 'h100217, 'h100218, 'h10003c, 'h100047, 'h10021a, 'h10021d, 'h10021b, 'h10021c, 'h10021e, 'h100221, 'h10021f, 'h2004f8, 'h100220, 'h1000b6, 'h100222, 'h100225, 'h1000b3, 'h1000b4, 'h100223, 'h1000b5, 'h100224, 'h1000b7, 'h100226, 'h100229, 'h10003c, 'h100047, 'h100227, 'h100228, 'h10022a, 'h10022d, 'h10022b, 'h10022c, 'h2004f8, 'h10022e, 'h100231, 'h10022f, 'h100230, 'h1000b6, 'h100232, 'h100235, 'h1000b3, 'h1000b4, 'h100233, 'h1000b5, 'h100234, 'h10003c, 'h100047, 'h1000b7, 'h100236, 'h100239, 'h100237, 'h100238, 'h10023a, 'h2004f8, 'h10023d, 'h10023b, 'h10023c, 'h10023e, 'h1000b6, 'h100241, 'h10023f, 'h1000b3, 'h1000b4, 'h100240, 'h1000b5, 'h100242, 'h10003c, 'h100047, 'h1000b7, 'h100246, 'h100243, 'h100244, 'h100245, 'h10024a, 'h2004f8, 'h100247, 'h100248, 'h100249, 'h10024e, 'h10024b, 'h10024c, 'h10024d, 'h1000b6, 'h100252, 'h1000b3, 'h10024f, 'h1000b4, 'h10003c, 'h100047, 'h100250, 'h1000b5, 'h100251, 'h1000b7, 'h100256, 'h100253, 'h2004f8, 'h100254, 'h100255, 'h10025a, 'h100257, 'h100258, 'h100259, 'h10025e, 'h10025b, 'h10025c, 'h10025d, 'h1000b6, 'h100262, 'h10003c, 'h100047, 'h1000b3, 'h10025f, 'h1000b4, 'h100260, 'h1000b5, 'h100261, 'h2004f8, 'h1000b7, 'h100266, 'h100263, 'h100264, 'h100265, 'h100267, 'h10026a, 'h100268, 'h100269, 'h10026b, 'h10026e, 'h10026c, 'h10003c, 'h100047, 'h10026d, 'h1000b6, 'h10026f, 'h100272, 'h1000b3, 'h1000b4, 'h2004f8, 'h100270, 'h1000b5, 'h100271, 'h1000b7, 'h100171, 'h1000bb, 'h100174, 'h1000b8, 'h100172, 'h1000b9, 'h100173, 'h1000ba, 'h10003c, 'h100047, 'h100175, 'h100178, 'h100176, 'h100177, 'h100179, 'h10017c, 'h2004f8, 'h10017a, 'h10017b, 'h10017d, 'h100180, 'h1000b7, 'h10017e, 'h10017f, 'h1000bb, 'h100181, 'h100184, 'h1000b8, 'h100182, 'h10003c, 'h100047, 'h1000b9, 'h100183, 'h1000ba, 'h100185, 'h100188, 'h100186, 'h2004f8, 'h100187, 'h100189, 'h10018c, 'h10018a, 'h10018b, 'h10018d, 'h100190, 'h1000bb, 'h1000b7, 'h10018e, 'h1000b8, 'h10018f, 'h10003c, 'h100047, 'h1000b9, 'h100191, 'h100194, 'h100192, 'h100193, 'h1000ba, 'h2004f8, 'h100195, 'h100198, 'h100196, 'h100197, 'h100199, 'h10019c, 'h10019a, 'h10019b, 'h1000bb, 'h10019d, 'h1001a0, 'h1000b7, 'h10003c, 'h100047, 'h1000b8, 'h10019e, 'h1000b9, 'h10019f, 'h1001a1, 'h1001a4, 'h2004f8, 'h1001a2, 'h1001a3, 'h1000ba, 'h1001a5, 'h1001a8, 'h1001a6, 'h1001a7, 'h1001a9, 'h1000bb, 'h1001ac, 'h1001aa, 'h1001ab, 'h10003c, 'h100047, 'h1001ad, 'h1001b0, 'h1000b7, 'h1000b8, 'h1001ae, 'h1000b9, 'h2004f8, 'h1001af, 'h1001b1, 'h1001b4, 'h1001b2, 'h1001b3, 'h1000ba, 'h1001b5, 'h1001b8, 'h1000bb, 'h1001b6, 'h1001b7, 'h1001b9, 'h10003c, 'h100047, 'h1001bc, 'h1001ba, 'h1001bb, 'h1001bd, 'h1001c1, 'h1000b7, 'h2004f8, 'h1001be, 'h1000b8, 'h1001bf, 'h1000b9, 'h1001c0, 'h1000ba, 'h1001c5, 'h1001c2, 'h1001c3, 'h1001c4, 'h1000bb, 'h1001c9, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001cd, 'h1001ca, 'h1000b7, 'h2004f8, 'h1001cb, 'h1000b8, 'h1001cc, 'h1000b9, 'h1001d1, 'h1001ce, 'h1001cf, 'h1001d0, 'h1000ba, 'h1001d5, 'h1000bb, 'h1001d2, 'h10003c, 'h100047, 'h1001d3, 'h1001d4, 'h1001d9, 'h1001d6, 'h1001d7, 'h1001d8, 'h2004f8, 'h1001dd, 'h1000b7, 'h1001da, 'h1000b8, 'h1001db, 'h1000b9, 'h1001dc, 'h1001e1, 'h1001de, 'h1001df, 'h1001e0, 'h1000ba, 'h10003c, 'h100047, 'h1000bb, 'h1001e2, 'h1001e5, 'h1001e3, 'h1001e4, 'h1001e6, 'h2004f8, 'h1001e9, 'h1000b7, 'h1001e7, 'h1000b8, 'h1001e8, 'h1000b9, 'h1001ea, 'h1001ed, 'h1001eb, 'h1001ec, 'h1001ee, 'h1001f1, 'h10003c, 'h100047, 'h1000bb, 'h1001ef, 'h1001f0, 'h1000ba, 'h1001f2, 'h1001f5, 'h2004f8, 'h1001f3, 'h1001f4, 'h1001f6, 'h1001f9, 'h1000b7, 'h1000b8, 'h1001f7, 'h1000b9, 'h1001f8, 'h1001fa, 'h1001fd, 'h1001fb, 'h10003c, 'h100047, 'h1001fc, 'h1000bb, 'h1001fe, 'h100201, 'h1001ff, 'h100200, 'h2004f8, 'h1000ba, 'h100202, 'h100205, 'h100203, 'h100204, 'h100206, 'h100209, 'h1000b7, 'h1000b8, 'h100207, 'h1000b9, 'h100208, 'h10003c, 'h100047, 'h10020a, 'h1000bb, 'h10020d, 'h10020b, 'h10020c, 'h10020e, 'h2004f8, 'h100211, 'h10020f, 'h100210, 'h1000ba, 'h100212, 'h100215, 'h100213, 'h100214, 'h100216, 'h100219, 'h1000b7, 'h1000b8, 'h10003c, 'h100047, 'h100217, 'h1000b9, 'h100218, 'h1000bb, 'h10021a, 'h10021d, 'h2004f8, 'h10021b, 'h10021c, 'h10021e, 'h100221, 'h10021f, 'h100220, 'h1000ba, 'h100222, 'h100225, 'h100223, 'h100224, 'h100226, 'h100229, 'h10003c, 'h100047, 'h1000b7, 'h1000b8, 'h100227, 'h1000b9, 'h100228, 'h2004f8, 'h1000bb, 'h10022a, 'h10022d, 'h10022b, 'h10022c, 'h10022e, 'h100231, 'h10022f, 'h100230, 'h1000ba, 'h100232, 'h100235, 'h100233, 'h10003c, 'h100047, 'h100234, 'h100236, 'h100239, 'h1000b7, 'h1000b8, 'h2004f8, 'h100237, 'h1000b9, 'h100238, 'h1000bb, 'h10023a, 'h10023d, 'h10023b, 'h10023c, 'h10023e, 'h100242, 'h10023f, 'h100240, 'h100241, 'h10003c, 'h100047, 'h1000ba, 'h100246, 'h100243, 'h1000b7, 'h1000b8, 'h2004f8, 'h100244, 'h1000b9, 'h100245, 'h1000bb, 'h10024a, 'h100247, 'h100248, 'h100249, 'h10024e, 'h10024b, 'h10024c, 'h10024d, 'h100252, 'h10003c, 'h100047, 'h10024f, 'h100250, 'h100251, 'h1000ba, 'h100256, 'h2004f8, 'h1000b7, 'h100253, 'h1000b8, 'h100254, 'h1000b9, 'h100255, 'h1000bb, 'h10025a, 'h100257, 'h100258, 'h100259, 'h10025e, 'h10025b, 'h10003c, 'h100047, 'h10025c, 'h10025d, 'h100262, 'h10025f, 'h100260, 'h2004f8, 'h100261, 'h1000ba, 'h100263, 'h100266, 'h1000b7, 'h1000b8, 'h100264, 'h1000b9, 'h100265, 'h1000bb, 'h100267, 'h10026a, 'h100268, 'h10003c, 'h100047, 'h100269, 'h10026b, 'h10026e, 'h10026c, 'h10026d, 'h2004f8, 'h10026f, 'h100272, 'h100270, 'h100271, 'h1000ba, 'h100171, 'h1000bf, 'h1000bc, 'h100172, 'h1000bd, 'h100173, 'h1000be, 'h100174, 'h10003c, 'h100047, 'h100175, 'h1000bb, 'h100176, 'h100177, 'h100178, 'h2004f8, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000bf, 'h100181, 'h1000bc, 'h100182, 'h1000bd, 'h10003c, 'h100047, 'h100183, 'h1000be, 'h100184, 'h100185, 'h1000bb, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h1000bf, 'h10018e, 'h1000bc, 'h10018f, 'h1000bd, 'h10003c, 'h100047, 'h100190, 'h1000be, 'h100191, 'h100192, 'h100193, 'h2004f8, 'h100194, 'h100195, 'h1000bb, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h1000bf, 'h10019d, 'h1000bc, 'h10003c, 'h100047, 'h10019e, 'h1000bd, 'h10019f, 'h1000be, 'h1001a0, 'h2004f8, 'h1001a1, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1000bb, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1000bf, 'h1001aa, 'h1000bc, 'h10003c, 'h100047, 'h1001ab, 'h1000bd, 'h1001ac, 'h1000be, 'h1001ad, 'h2004f8, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1000bb, 'h1001b6, 'h1001b7, 'h1001b8, 'h1000bf, 'h10003c, 'h100047, 'h1001b9, 'h1000bc, 'h1001ba, 'h1000bd, 'h1001bb, 'h2004f8, 'h1000be, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1000bb, 'h1001c3, 'h1001c4, 'h1001c5, 'h1000bf, 'h10003c, 'h100047, 'h1001c6, 'h1000bc, 'h1001c7, 'h1000bd, 'h1001c8, 'h2004f8, 'h1000be, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1000bb, 'h1001d2, 'h1001d3, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1000bf, 'h1001d6, 'h1000bc, 'h2004f8, 'h1001d7, 'h1000bd, 'h1001d8, 'h1000be, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1000bb, 'h1001df, 'h1001e0, 'h10003c, 'h100047, 'h1001e1, 'h1001e2, 'h1000bf, 'h1001e3, 'h1000bc, 'h2004f8, 'h1001e4, 'h1000bd, 'h1001e5, 'h1000be, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h10003c, 'h100047, 'h1000bb, 'h1001ef, 'h1001f0, 'h1001f1, 'h1000bf, 'h2004f8, 'h1001f2, 'h1000bc, 'h1001f3, 'h1000bd, 'h1001f4, 'h1000be, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h10003c, 'h100047, 'h1001fc, 'h1001fd, 'h1001fe, 'h1000bb, 'h1001ff, 'h2004f8, 'h100200, 'h100201, 'h1000bf, 'h100202, 'h1000bc, 'h100203, 'h1000bd, 'h100204, 'h1000be, 'h100205, 'h100206, 'h100207, 'h100208, 'h10003c, 'h100047, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h2004f8, 'h10020e, 'h1000bb, 'h10020f, 'h100210, 'h100211, 'h1000bf, 'h100212, 'h1000bc, 'h100213, 'h1000bd, 'h100214, 'h1000be, 'h100215, 'h10003c, 'h100047, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h2004f8, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h1000bb, 'h10021f, 'h100220, 'h100221, 'h1000bf, 'h100222, 'h1000bc, 'h100223, 'h1000bd, 'h10003c, 'h100047, 'h100224, 'h1000be, 'h100225, 'h100226, 'h100227, 'h2004f8, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h1000bb, 'h10022f, 'h100230, 'h100231, 'h1000bf, 'h100232, 'h10003c, 'h100047, 'h1000bc, 'h100233, 'h1000bd, 'h100234, 'h1000be, 'h2004f8, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h1000bb, 'h10023f, 'h100240, 'h10003c, 'h100047, 'h100241, 'h100242, 'h1000bf, 'h100243, 'h1000bc, 'h2004f8, 'h100244, 'h1000bd, 'h100245, 'h1000be, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h1000bb, 'h10024c, 'h10024d, 'h10003c, 'h100047, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h2004f8, 'h1000bf, 'h100253, 'h1000bc, 'h100254, 'h1000bd, 'h100255, 'h1000be, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h1000bb, 'h10003c, 'h100047, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h2004f8, 'h1000bf, 'h100260, 'h1000bc, 'h100261, 'h1000bd, 'h100262, 'h1000be, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10003c, 'h100047, 'h10026a, 'h10026b, 'h1000bb, 'h10026c, 'h2004f8, 'h10026d, 'h10026e, 'h1000bf, 'h10026f, 'h1000bc, 'h100270, 'h1000bd, 'h100271, 'h1000be, 'h100272, 'h100171, 'h1000c3, 'h100173, 'h1000c0, 'h10003c, 'h100047, 'h100172, 'h1000c1, 'h1000c2, 'h100174, 'h2004f8, 'h100175, 'h100177, 'h1000bf, 'h100176, 'h100178, 'h100179, 'h10017b, 'h10017a, 'h10017c, 'h10017d, 'h10017f, 'h1000c3, 'h10017e, 'h1000c0, 'h10003c, 'h100047, 'h100180, 'h100181, 'h100183, 'h100182, 'h2004f8, 'h1000c1, 'h1000c2, 'h100184, 'h100185, 'h100187, 'h1000bf, 'h100186, 'h100188, 'h100189, 'h10018b, 'h10018a, 'h10018c, 'h1000c3, 'h10018d, 'h10018f, 'h10003c, 'h100047, 'h1000c0, 'h10018e, 'h100190, 'h2004f8, 'h100191, 'h100193, 'h100192, 'h1000c1, 'h1000c2, 'h100194, 'h100195, 'h100197, 'h1000bf, 'h100196, 'h100198, 'h100199, 'h1000c3, 'h10019c, 'h10019a, 'h10003c, 'h100047, 'h1000c0, 'h10019b, 'h10019d, 'h2004f8, 'h1001a0, 'h10019e, 'h10019f, 'h1000c1, 'h1000c2, 'h1001a1, 'h1001a4, 'h1001a2, 'h1001a3, 'h1001a5, 'h1001a8, 'h1000bf, 'h1001a6, 'h1001a7, 'h1000c3, 'h10003c, 'h100047, 'h1001a9, 'h1001ac, 'h1000c0, 'h2004f8, 'h1001aa, 'h1001ab, 'h1001ad, 'h1001b0, 'h1001ae, 'h1000c1, 'h1001af, 'h1000c2, 'h1001b1, 'h1001b4, 'h1001b2, 'h1001b3, 'h1001b5, 'h1001b8, 'h1000c3, 'h10003c, 'h100047, 'h1000bf, 'h1001b6, 'h1000c0, 'h2004f8, 'h1001b7, 'h1001b9, 'h1001bc, 'h1001ba, 'h1001bb, 'h1000c1, 'h1001bd, 'h1001c0, 'h1001be, 'h1001bf, 'h1000c2, 'h1001c1, 'h1001c4, 'h1001c2, 'h1001c3, 'h10003c, 'h100047, 'h1001c5, 'h1000c3, 'h1001c8, 'h2004f8, 'h1000bf, 'h1001c6, 'h1000c0, 'h1001c7, 'h1001c9, 'h1001cc, 'h1001ca, 'h1001cb, 'h1000c1, 'h1001cd, 'h1000c2, 'h1001d0, 'h1001ce, 'h1001cf, 'h1001d1, 'h10003c, 'h100047, 'h1001d4, 'h1000c3, 'h1001d2, 'h2004f8, 'h1000bf, 'h1001d3, 'h1000c0, 'h1001d5, 'h1001d8, 'h1001d6, 'h1001d7, 'h1001d9, 'h1001da, 'h1001dc, 'h1001db, 'h1000c1, 'h1000c2, 'h1001dd, 'h1001de, 'h1001e0, 'h10003c, 'h100047, 'h1000c3, 'h1001df, 'h2004f8, 'h1001e1, 'h1001e2, 'h1001e4, 'h1000bf, 'h1000c0, 'h1001e3, 'h1001e5, 'h1001e6, 'h1001e8, 'h1001e7, 'h1001e9, 'h1001ea, 'h1001ec, 'h1001eb, 'h1000c1, 'h1000c2, 'h10003c, 'h100047, 'h1001ed, 'h1000c3, 'h2004f8, 'h1001ee, 'h1001f0, 'h1001ef, 'h1001f1, 'h1001f2, 'h1001f4, 'h1000bf, 'h1000c0, 'h1001f3, 'h1001f5, 'h1001f6, 'h1001f8, 'h1001f7, 'h1001f9, 'h1001fa, 'h1001fc, 'h10003c, 'h100047, 'h1001fb, 'h1000c1, 'h2004f8, 'h1000c2, 'h1001fd, 'h1000c3, 'h1001fe, 'h100200, 'h1001ff, 'h100201, 'h100202, 'h100204, 'h1000bf, 'h1000c0, 'h100203, 'h100205, 'h100206, 'h100208, 'h100207, 'h10003c, 'h100047, 'h100209, 'h10020a, 'h2004f8, 'h10020c, 'h10020b, 'h1000c1, 'h1000c2, 'h10020d, 'h1000c3, 'h10020e, 'h100210, 'h10020f, 'h100211, 'h100212, 'h100214, 'h1000bf, 'h1000c0, 'h100213, 'h100215, 'h10003c, 'h100047, 'h100216, 'h100218, 'h2004f8, 'h100217, 'h100219, 'h10021a, 'h10021d, 'h10021b, 'h1000c1, 'h10021c, 'h1000c2, 'h1000c3, 'h10021e, 'h100221, 'h10021f, 'h100220, 'h100222, 'h100225, 'h1000bf, 'h10003c, 'h100047, 'h1000c0, 'h100223, 'h2004f8, 'h100224, 'h100226, 'h100229, 'h100227, 'h100228, 'h1000c1, 'h10022a, 'h10022d, 'h1000c3, 'h10022b, 'h10022c, 'h1000c2, 'h10022e, 'h100231, 'h10022f, 'h100230, 'h10003c, 'h100047, 'h100232, 'h100235, 'h2004f8, 'h1000bf, 'h1000c0, 'h100233, 'h100234, 'h100236, 'h100239, 'h100237, 'h1000c1, 'h100238, 'h1000c3, 'h10023a, 'h10023d, 'h10023b, 'h10023c, 'h1000c2, 'h10023e, 'h10003c, 'h100047, 'h100241, 'h10023f, 'h2004f8, 'h100240, 'h100242, 'h100245, 'h1000bf, 'h100243, 'h1000c0, 'h100244, 'h1000c1, 'h100246, 'h1000c3, 'h100249, 'h100247, 'h100248, 'h10024a, 'h1000c2, 'h10024d, 'h10003c, 'h100047, 'h10024b, 'h10024c, 'h2004f8, 'h10024e, 'h100251, 'h10024f, 'h1000bf, 'h100250, 'h1000c0, 'h100252, 'h100255, 'h100253, 'h100254, 'h1000c1, 'h100256, 'h1000c3, 'h100259, 'h100257, 'h100258, 'h10003c, 'h100047, 'h1000c2, 'h10025a, 'h2004f8, 'h10025b, 'h10025d, 'h10025c, 'h10025e, 'h10025f, 'h100261, 'h1000bf, 'h1000c0, 'h100260, 'h100262, 'h100263, 'h100265, 'h1000c3, 'h100264, 'h1000c1, 'h100266, 'h10003c, 'h100047, 'h1000c2, 'h100267, 'h2004f8, 'h100269, 'h100268, 'h10026a, 'h10026b, 'h10026d, 'h10026c, 'h10026e, 'h10026f, 'h100271, 'h1000bf, 'h1000c0, 'h100270, 'h100272, 'h1000c3, 'h100171, 'h1000c7, 'h10003c, 'h100047, 'h1000c4, 'h100172, 'h2004f8, 'h1000c5, 'h100173, 'h1000c6, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h1000c3, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h100180, 'h1000c7, 'h2004f8, 'h100181, 'h1000c4, 'h100182, 'h1000c5, 'h100183, 'h1000c6, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h1000c3, 'h10018e, 'h2004f8, 'h10018f, 'h100190, 'h1000c7, 'h100191, 'h1000c4, 'h100192, 'h1000c5, 'h100193, 'h1000c6, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10003c, 'h100047, 'h10019b, 'h10019c, 'h2004f8, 'h10019d, 'h1000c3, 'h10019e, 'h10019f, 'h1001a0, 'h1000c7, 'h1001a1, 'h1000c4, 'h1001a2, 'h1000c5, 'h1001a3, 'h1000c6, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h10003c, 'h100047, 'h1001a8, 'h1001a9, 'h2004f8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1000c3, 'h1001ae, 'h1001af, 'h1001b0, 'h1000c7, 'h1001b1, 'h1000c4, 'h1001b2, 'h1000c5, 'h1001b3, 'h1000c6, 'h1001b4, 'h10003c, 'h100047, 'h1001b5, 'h1001b6, 'h2004f8, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1000c3, 'h1001be, 'h1001bf, 'h1001c0, 'h1000c7, 'h1001c1, 'h1000c4, 'h1001c2, 'h1000c5, 'h10003c, 'h100047, 'h1001c3, 'h1000c6, 'h2004f8, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1000c3, 'h1001cb, 'h1001cc, 'h1001cd, 'h1000c7, 'h1001ce, 'h1000c4, 'h1001cf, 'h1000c5, 'h10003c, 'h100047, 'h1001d0, 'h1000c6, 'h2004f8, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1000c3, 'h1001db, 'h1001dc, 'h1001dd, 'h1000c7, 'h1001de, 'h10003c, 'h100047, 'h1000c4, 'h1001df, 'h2004f8, 'h1000c5, 'h1001e0, 'h1000c6, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1000c3, 'h1001eb, 'h1001ec, 'h10003c, 'h100047, 'h1001ed, 'h1000c7, 'h2004f8, 'h1001ee, 'h1000c4, 'h1001ef, 'h1000c5, 'h1001f0, 'h1000c6, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h10003c, 'h100047, 'h1000c3, 'h1001fb, 'h2004f8, 'h1001fc, 'h1001fd, 'h1000c7, 'h1001fe, 'h1000c4, 'h1001ff, 'h1000c5, 'h100200, 'h1000c6, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100207, 'h10003c, 'h100047, 'h100208, 'h100209, 'h2004f8, 'h10020a, 'h1000c3, 'h10020b, 'h10020c, 'h10020d, 'h1000c7, 'h10020e, 'h1000c4, 'h10020f, 'h1000c5, 'h100210, 'h1000c6, 'h100211, 'h100212, 'h100213, 'h100214, 'h10003c, 'h100047, 'h100215, 'h100216, 'h2004f8, 'h100217, 'h100218, 'h100219, 'h10021a, 'h1000c3, 'h10021b, 'h10021c, 'h10021d, 'h1000c7, 'h10021e, 'h1000c4, 'h10021f, 'h1000c5, 'h100220, 'h1000c6, 'h100221, 'h10003c, 'h100047, 'h100222, 'h100223, 'h2004f8, 'h100224, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h1000c3, 'h10022b, 'h10022c, 'h10022d, 'h1000c7, 'h10022e, 'h1000c4, 'h10022f, 'h1000c5, 'h10003c, 'h100047, 'h100230, 'h1000c6, 'h2004f8, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h1000c3, 'h10023b, 'h10023c, 'h10023d, 'h1000c7, 'h10023e, 'h10003c, 'h100047, 'h1000c4, 'h10023f, 'h2004f8, 'h1000c5, 'h100240, 'h1000c6, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h1000c3, 'h10024b, 'h10024c, 'h10003c, 'h100047, 'h10024d, 'h10024e, 'h2004f8, 'h1000c7, 'h10024f, 'h1000c4, 'h100250, 'h1000c5, 'h100251, 'h1000c6, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h1000c3, 'h100258, 'h100259, 'h10003c, 'h100047, 'h10025a, 'h10025b, 'h2004f8, 'h1000c7, 'h10025c, 'h1000c4, 'h10025d, 'h1000c5, 'h10025e, 'h1000c6, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h10003c, 'h100047, 'h1000c3, 'h100268, 'h2004f8, 'h100269, 'h10026a, 'h1000c7, 'h10026b, 'h1000c4, 'h10026c, 'h1000c5, 'h10026d, 'h1000c6, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000cb, 'h10003c, 'h100047, 'h1000c8, 'h100172, 'h2004f8, 'h1000c9, 'h100173, 'h1000ca, 'h100174, 'h100175, 'h1000c7, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h100180, 'h1000cb, 'h2004f8, 'h100181, 'h1000c8, 'h100182, 'h1000c9, 'h100183, 'h1000ca, 'h100184, 'h100185, 'h1000c7, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10003c, 'h100047, 'h10018d, 'h1000cb, 'h2004f8, 'h10018e, 'h1000c8, 'h10018f, 'h1000c9, 'h100190, 'h1000ca, 'h100191, 'h100192, 'h100193, 'h100194, 'h100195, 'h1000c7, 'h100196, 'h100197, 'h100198, 'h100199, 'h10003c, 'h100047, 'h10019a, 'h10019b, 'h2004f8, 'h10019c, 'h1000cb, 'h10019d, 'h1000c8, 'h10019e, 'h1000c9, 'h10019f, 'h1000ca, 'h1001a0, 'h1001a1, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1000c7, 'h1001a6, 'h10003c, 'h100047, 'h1001a7, 'h1001a8, 'h2004f8, 'h1001a9, 'h1000cb, 'h1001aa, 'h1000c8, 'h1001ab, 'h1000c9, 'h1001ac, 'h1000ca, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h10003c, 'h100047, 'h1001b5, 'h1000c7, 'h2004f8, 'h1001b6, 'h1001b7, 'h1001b8, 'h1000cb, 'h1001b9, 'h1000c8, 'h1001ba, 'h1000c9, 'h1001bb, 'h1000ca, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h10003c, 'h100047, 'h1001c2, 'h1001c3, 'h2004f8, 'h1001c4, 'h1001c5, 'h1000c7, 'h1001c6, 'h1001c7, 'h1001c8, 'h1000cb, 'h1001c9, 'h1001ca, 'h1000c8, 'h1001cb, 'h1000c9, 'h1001cc, 'h1000ca, 'h1001cd, 'h1001ce, 'h10003c, 'h100047, 'h1001cf, 'h1001d0, 'h2004f8, 'h1001d1, 'h1001d2, 'h1000c7, 'h1001d3, 'h1001d4, 'h1001d5, 'h1000cb, 'h1001d6, 'h1001d7, 'h1000c8, 'h1001d8, 'h1000c9, 'h1001d9, 'h1000ca, 'h1001da, 'h1001db, 'h10003c, 'h100047, 'h1001dc, 'h1001dd, 'h2004f8, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000c7, 'h1001e3, 'h1001e4, 'h1001e5, 'h1000cb, 'h1001e6, 'h1000c8, 'h1001e7, 'h1000c9, 'h1001e8, 'h1000ca, 'h10003c, 'h100047, 'h1001e9, 'h1001ea, 'h2004f8, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000c7, 'h1001f3, 'h1001f4, 'h1001f5, 'h1000cb, 'h1001f6, 'h1000c8, 'h1001f7, 'h10003c, 'h100047, 'h1000c9, 'h1001f8, 'h2004f8, 'h1000ca, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h1000c7, 'h100203, 'h100204, 'h100205, 'h1000cb, 'h10003c, 'h100047, 'h100206, 'h1000c8, 'h2004f8, 'h100207, 'h1000c9, 'h100208, 'h1000ca, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000c7, 'h100213, 'h10003c, 'h100047, 'h100214, 'h100215, 'h2004f8, 'h1000cb, 'h100216, 'h1000c8, 'h100217, 'h1000c9, 'h100218, 'h1000ca, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h10003c, 'h100047, 'h100222, 'h1000c7, 'h2004f8, 'h100223, 'h100224, 'h100225, 'h1000cb, 'h100226, 'h1000c8, 'h100227, 'h1000c9, 'h100228, 'h1000ca, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10003c, 'h100047, 'h10022f, 'h100230, 'h2004f8, 'h100231, 'h100232, 'h1000c7, 'h100233, 'h100234, 'h100235, 'h1000cb, 'h100236, 'h1000c8, 'h100237, 'h1000c9, 'h100238, 'h1000ca, 'h100239, 'h10023a, 'h10023b, 'h10003c, 'h100047, 'h10023c, 'h10023d, 'h2004f8, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h1000c7, 'h100243, 'h100244, 'h100245, 'h1000cb, 'h100246, 'h1000c8, 'h100247, 'h1000c9, 'h100248, 'h1000ca, 'h10003c, 'h100047, 'h100249, 'h10024a, 'h2004f8, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h1000c7, 'h100250, 'h100251, 'h100252, 'h1000cb, 'h100253, 'h1000c8, 'h100254, 'h1000c9, 'h100255, 'h1000ca, 'h10003c, 'h100047, 'h100256, 'h100257, 'h2004f8, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h1000c7, 'h100260, 'h100261, 'h100262, 'h1000cb, 'h100263, 'h1000c8, 'h100264, 'h10003c, 'h100047, 'h1000c9, 'h100265, 'h2004f8, 'h1000ca, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h1000c7, 'h100270, 'h100271, 'h100272, 'h1000cb, 'h10003c, 'h100047, 'h100171, 'h1000cf, 'h2004f8, 'h1000cc, 'h100172, 'h1000cd, 'h100173, 'h1000ce, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10003c, 'h100047, 'h10017f, 'h100180, 'h2004f8, 'h1000cf, 'h100181, 'h1000cc, 'h100182, 'h1000cd, 'h100183, 'h1000ce, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10003c, 'h100047, 'h10018d, 'h10018e, 'h2004f8, 'h10018f, 'h100190, 'h1000cf, 'h100191, 'h1000cc, 'h100192, 'h1000cd, 'h100193, 'h1000ce, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10003c, 'h100047, 'h10019b, 'h10019c, 'h2004f8, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1000cf, 'h1001a1, 'h1000cc, 'h1001a2, 'h1000cd, 'h1001a3, 'h1000ce, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h10003c, 'h100047, 'h1001a9, 'h1001aa, 'h2004f8, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1000cf, 'h1001b1, 'h1000cc, 'h1001b2, 'h1000cd, 'h1001b3, 'h1000ce, 'h1001b4, 'h1001b5, 'h1001b6, 'h10003c, 'h100047, 'h1001b7, 'h1001b8, 'h2004f8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1000cf, 'h1001c1, 'h1000cc, 'h1001c2, 'h1000cd, 'h1001c3, 'h1000ce, 'h1001c4, 'h10003c, 'h100047, 'h1001c5, 'h1001c6, 'h2004f8, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1000cf, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000cc, 'h1001d3, 'h1000cd, 'h10003c, 'h100047, 'h1001d4, 'h1000ce, 'h2004f8, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1000cf, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000cc, 'h10003c, 'h100047, 'h1001e3, 'h1000cd, 'h2004f8, 'h1001e4, 'h1000ce, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1000cf, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h10003c, 'h100047, 'h1001f2, 'h1000cc, 'h2004f8, 'h1001f3, 'h1000cd, 'h1001f4, 'h1000ce, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1000cf, 'h1001fe, 'h1001ff, 'h10003c, 'h100047, 'h100200, 'h100201, 'h2004f8, 'h100202, 'h1000cc, 'h100203, 'h1000cd, 'h100204, 'h1000ce, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h1000cf, 'h10003c, 'h100047, 'h10020e, 'h10020f, 'h2004f8, 'h100210, 'h100211, 'h100212, 'h1000cc, 'h100213, 'h1000cd, 'h100214, 'h1000ce, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10003c, 'h100047, 'h10021d, 'h1000cf, 'h2004f8, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000cc, 'h100223, 'h1000cd, 'h100224, 'h1000ce, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10003c, 'h100047, 'h10022b, 'h10022c, 'h2004f8, 'h10022d, 'h1000cf, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h1000cc, 'h100233, 'h1000cd, 'h100234, 'h1000ce, 'h100235, 'h100236, 'h100237, 'h100238, 'h10003c, 'h100047, 'h100239, 'h10023a, 'h2004f8, 'h10023b, 'h10023c, 'h10023d, 'h1000cf, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h1000cc, 'h100243, 'h1000cd, 'h100244, 'h1000ce, 'h100245, 'h100246, 'h10003c, 'h100047, 'h100247, 'h100248, 'h2004f8, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h1000cf, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h1000cc, 'h100254, 'h1000cd, 'h100255, 'h10003c, 'h100047, 'h1000ce, 'h100256, 'h2004f8, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h1000cf, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h1000cc, 'h100264, 'h10003c, 'h100047, 'h1000cd, 'h100265, 'h2004f8, 'h1000ce, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h1000cf, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000d3, 'h10003c, 'h100047, 'h1000d0, 'h2004f8, 'h100172, 'h1000d1, 'h100173, 'h1000d2, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h10003c, 'h100047, 'h1000d3, 'h2004f8, 'h100181, 'h1000d0, 'h100182, 'h1000d1, 'h100183, 'h1000d2, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10003c, 'h100047, 'h10018f, 'h2004f8, 'h100190, 'h1000d3, 'h100191, 'h1000d0, 'h100192, 'h1000d1, 'h100193, 'h1000d2, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10003c, 'h100047, 'h10019d, 'h2004f8, 'h10019e, 'h10019f, 'h1001a0, 'h1000d3, 'h1001a1, 'h1000d0, 'h1001a2, 'h1000d1, 'h1001a3, 'h1000d2, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h10003c, 'h100047, 'h1001ab, 'h2004f8, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1000d3, 'h1001b1, 'h1000d0, 'h1001b2, 'h1000d1, 'h1001b3, 'h1000d2, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h10003c, 'h100047, 'h1001b9, 'h2004f8, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1000d3, 'h1001c1, 'h1000d0, 'h1001c2, 'h1000d1, 'h1001c3, 'h1000d2, 'h1001c4, 'h1001c5, 'h1001c6, 'h10003c, 'h100047, 'h1001c7, 'h2004f8, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1000d3, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000d0, 'h1001d3, 'h1000d1, 'h1001d4, 'h1000d2, 'h10003c, 'h100047, 'h1001d5, 'h2004f8, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1000d3, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000d0, 'h1001e3, 'h1000d1, 'h10003c, 'h100047, 'h1001e4, 'h2004f8, 'h1000d2, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1000d3, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000d0, 'h10003c, 'h100047, 'h1001f3, 'h2004f8, 'h1000d1, 'h1001f4, 'h1000d2, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1000d3, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h10003c, 'h100047, 'h100202, 'h2004f8, 'h1000d0, 'h100203, 'h1000d1, 'h100204, 'h1000d2, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h1000d3, 'h10020e, 'h10020f, 'h10003c, 'h100047, 'h100210, 'h2004f8, 'h100211, 'h100212, 'h1000d0, 'h100213, 'h1000d1, 'h100214, 'h1000d2, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h1000d3, 'h10003c, 'h100047, 'h10021e, 'h2004f8, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000d0, 'h100223, 'h1000d1, 'h100224, 'h1000d2, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10003c, 'h100047, 'h10022d, 'h2004f8, 'h1000d3, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h1000d0, 'h100233, 'h1000d1, 'h100234, 'h1000d2, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10003c, 'h100047, 'h10023b, 'h2004f8, 'h10023c, 'h10023d, 'h1000d3, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h1000d0, 'h100243, 'h1000d1, 'h100244, 'h1000d2, 'h100245, 'h100246, 'h100247, 'h100248, 'h10003c, 'h100047, 'h100249, 'h2004f8, 'h10024a, 'h10024b, 'h1000d3, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h1000d0, 'h100254, 'h1000d1, 'h100255, 'h1000d2, 'h100256, 'h10003c, 'h100047, 'h100257, 'h2004f8, 'h100258, 'h100259, 'h10025a, 'h1000d3, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h1000d0, 'h100264, 'h1000d1, 'h100265, 'h10003c, 'h100047, 'h1000d2, 'h2004f8, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h1000d3, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000d7, 'h1000d4, 'h10003c, 'h100047, 'h100172, 'h2004f8, 'h1000d5, 'h100173, 'h1000d6, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000d7, 'h10003c, 'h100047, 'h100181, 'h2004f8, 'h1000d4, 'h100182, 'h1000d5, 'h100183, 'h1000d6, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h10003c, 'h100047, 'h100190, 'h2004f8, 'h1000d7, 'h100191, 'h1000d4, 'h100192, 'h1000d5, 'h100193, 'h1000d6, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10003c, 'h100047, 'h10019e, 'h2004f8, 'h10019f, 'h1001a0, 'h1000d7, 'h1001a1, 'h1000d4, 'h1001a2, 'h1000d5, 'h1001a3, 'h1000d6, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h10003c, 'h100047, 'h1001ac, 'h2004f8, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1000d7, 'h1001b1, 'h1000d4, 'h1001b2, 'h1000d5, 'h1001b3, 'h1000d6, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h10003c, 'h100047, 'h1001ba, 'h2004f8, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1000d7, 'h1001c1, 'h1001c2, 'h1000d4, 'h1000d5, 'h1001c3, 'h1000d6, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h10003c, 'h100047, 'h1001c8, 'h2004f8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1000d7, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000d4, 'h1000d5, 'h1001d3, 'h1000d6, 'h1001d4, 'h1001d5, 'h10003c, 'h100047, 'h1001d6, 'h2004f8, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1000d7, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000d4, 'h1001e3, 'h1000d5, 'h1001e4, 'h10003c, 'h100047, 'h1000d6, 'h2004f8, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1000d7, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000d4, 'h1001f3, 'h10003c, 'h100047, 'h1000d5, 'h2004f8, 'h1001f4, 'h1000d6, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1000d7, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h10003c, 'h100047, 'h1000d4, 'h2004f8, 'h100203, 'h1000d5, 'h100204, 'h1000d6, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h1000d7, 'h10020e, 'h10020f, 'h100210, 'h10003c, 'h100047, 'h100211, 'h2004f8, 'h100212, 'h1000d4, 'h100213, 'h1000d5, 'h100214, 'h1000d6, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h1000d7, 'h10021e, 'h10003c, 'h100047, 'h10021f, 'h2004f8, 'h100220, 'h100221, 'h100222, 'h1000d4, 'h100223, 'h1000d5, 'h100224, 'h1000d6, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10003c, 'h100047, 'h1000d7, 'h2004f8, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h1000d4, 'h100233, 'h1000d5, 'h100234, 'h1000d6, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10003c, 'h100047, 'h10023c, 'h2004f8, 'h10023d, 'h1000d7, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h1000d4, 'h1000d5, 'h100244, 'h1000d6, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10003c, 'h100047, 'h10024a, 'h2004f8, 'h10024b, 'h1000d7, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h1000d4, 'h1000d5, 'h100254, 'h1000d6, 'h100255, 'h100256, 'h100257, 'h10003c, 'h100047, 'h100258, 'h2004f8, 'h100259, 'h10025a, 'h1000d7, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h1000d4, 'h100264, 'h1000d5, 'h100265, 'h1000d6, 'h10003c, 'h100047, 'h100266, 'h2004f8, 'h100267, 'h100268, 'h100269, 'h10026a, 'h1000d7, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000db, 'h1000d8, 'h100172, 'h10003c, 'h100047, 'h1000d9, 'h2004f8, 'h100173, 'h1000da, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000db, 'h100181, 'h10003c, 'h100047, 'h1000d8, 'h2004f8, 'h100182, 'h1000d9, 'h100183, 'h1000da, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h100190, 'h10003c, 'h100047, 'h1000db, 'h2004f8, 'h100191, 'h1000d8, 'h100192, 'h1000d9, 'h100193, 'h1000da, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10019e, 'h10003c, 'h100047, 'h10019f, 'h2004f8, 'h1001a0, 'h1000db, 'h1001a1, 'h1000d8, 'h1001a2, 'h1000d9, 'h1001a3, 'h1000da, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h10003c, 'h100047, 'h1001ad, 'h2004f8, 'h1001ae, 'h1001af, 'h1001b0, 'h1000db, 'h1001b1, 'h1000d8, 'h1001b2, 'h1000d9, 'h1001b3, 'h1000da, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h10003c, 'h100047, 'h1001bb, 'h2004f8, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1000db, 'h1001c1, 'h1001c2, 'h1000d8, 'h1000d9, 'h1001c3, 'h1000da, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h10003c, 'h100047, 'h1001c9, 'h2004f8, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1000db, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000d8, 'h1000d9, 'h1001d3, 'h1000da, 'h1001d4, 'h1001d5, 'h1001d6, 'h10003c, 'h100047, 'h1001d7, 'h2004f8, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1000db, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000d8, 'h1001e3, 'h1000d9, 'h1001e4, 'h1000da, 'h10003c, 'h100047, 'h1001e5, 'h2004f8, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1000db, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000d8, 'h1001f3, 'h1000d9, 'h10003c, 'h100047, 'h1001f4, 'h2004f8, 'h1000da, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1000db, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h1000d8, 'h10003c, 'h100047, 'h100203, 'h2004f8, 'h1000d9, 'h100204, 'h1000da, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h1000db, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h10003c, 'h100047, 'h100212, 'h2004f8, 'h1000d8, 'h100213, 'h1000d9, 'h100214, 'h1000da, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h1000db, 'h10021e, 'h10021f, 'h10003c, 'h100047, 'h100220, 'h2004f8, 'h100221, 'h100222, 'h1000d8, 'h100223, 'h1000d9, 'h100224, 'h1000da, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h1000db, 'h10003c, 'h100047, 'h10022e, 'h2004f8, 'h10022f, 'h100230, 'h100231, 'h100232, 'h1000d8, 'h100233, 'h1000d9, 'h100234, 'h1000da, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10003c, 'h100047, 'h10023d, 'h2004f8, 'h1000db, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h1000d8, 'h1000d9, 'h100244, 'h1000da, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10003c, 'h100047, 'h10024b, 'h2004f8, 'h1000db, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h1000d8, 'h1000d9, 'h100254, 'h1000da, 'h100255, 'h100256, 'h100257, 'h100258, 'h10003c, 'h100047, 'h100259, 'h2004f8, 'h1000db, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h1000d8, 'h100264, 'h1000d9, 'h100265, 'h1000da, 'h100266, 'h10003c, 'h100047, 'h100267, 'h2004f8, 'h1000db, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000df, 'h100172, 'h1000dc, 'h1000dd, 'h10003c, 'h100047, 'h100173, 'h2004f8, 'h1000de, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000df, 'h100181, 'h100182, 'h10003c, 'h100047, 'h1000dc, 'h2004f8, 'h1000dd, 'h100183, 'h1000de, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h1000df, 'h10018f, 'h100190, 'h10003c, 'h100047, 'h100191, 'h2004f8, 'h100192, 'h1000dc, 'h1000dd, 'h100193, 'h1000de, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h1000df, 'h10019d, 'h10019e, 'h10003c, 'h100047, 'h10019f, 'h2004f8, 'h1001a0, 'h1001a1, 'h1001a2, 'h1000dc, 'h1000dd, 'h1001a3, 'h1000de, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001ab, 'h1000df, 'h1001aa, 'h1001ac, 'h10003c, 'h100047, 'h1001ad, 'h2004f8, 'h1001af, 'h1001ae, 'h1001b0, 'h1001b1, 'h1001b3, 'h1000dc, 'h1001b2, 'h1000dd, 'h1000de, 'h1001b4, 'h1001b5, 'h1001b7, 'h1001b6, 'h1001b8, 'h1000df, 'h1001b9, 'h1001bb, 'h10003c, 'h100047, 'h1001ba, 'h2004f8, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1000dc, 'h1000dd, 'h1000de, 'h1001c4, 'h1001c5, 'h1001c6, 'h1000df, 'h1001c7, 'h1001c8, 'h10003c, 'h100047, 'h1001c9, 'h2004f8, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1000dc, 'h1000dd, 'h1000de, 'h1001d4, 'h1000df, 'h1001d5, 'h1001d6, 'h1001d7, 'h10003c, 'h100047, 'h2004f8, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1000dc, 'h1000dd, 'h1001e4, 'h1000de, 'h1001e5, 'h1000df, 'h10003c, 'h100047, 'h2004f8, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1000dc, 'h1000dd, 'h1001f4, 'h1000de, 'h10003c, 'h100047, 'h2004f8, 'h1001f5, 'h1000df, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h1000dc, 'h1000dd, 'h10003c, 'h100047, 'h2004f8, 'h100204, 'h1000de, 'h100205, 'h1000df, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100213, 'h10003c, 'h100047, 'h2004f8, 'h1000dc, 'h1000dd, 'h100214, 'h1000de, 'h100215, 'h1000df, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h10003c, 'h100047, 'h2004f8, 'h100222, 'h100223, 'h1000dc, 'h1000dd, 'h100224, 'h1000de, 'h100225, 'h1000df, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022c, 'h10022b, 'h10022d, 'h10022e, 'h100230, 'h10003c, 'h100047, 'h2004f8, 'h10022f, 'h100231, 'h100232, 'h100234, 'h1000dc, 'h100233, 'h1000dd, 'h1000de, 'h100235, 'h1000df, 'h100236, 'h100238, 'h100237, 'h100239, 'h10023a, 'h10023c, 'h10023b, 'h10023d, 'h10003c, 'h100047, 'h2004f8, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h1000dc, 'h1000dd, 'h1000de, 'h100245, 'h1000df, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10003c, 'h2004f8, 'h100047, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h1000dc, 'h1000dd, 'h1000de, 'h100255, 'h1000df, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10003c, 'h2004f8, 'h100047, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h1000dc, 'h1000dd, 'h100265, 'h1000de, 'h100266, 'h1000df, 'h100267, 'h100268, 'h10003c, 'h2004f8, 'h100047, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000e3, 'h1000e0, 'h100172, 'h1000e1, 'h100173, 'h1000e2, 'h100174, 'h10003c, 'h2004f8, 'h100047, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000e3, 'h100181, 'h1000e0, 'h100182, 'h1000e1, 'h100183, 'h10003c, 'h2004f8, 'h100047, 'h1000e2, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h100190, 'h1000e3, 'h100191, 'h1000e0, 'h100192, 'h10003c, 'h2004f8, 'h100047, 'h1000e1, 'h100193, 'h1000e2, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1000e3, 'h1001a1, 'h10003c, 'h2004f8, 'h100047, 'h1000e0, 'h1001a2, 'h1000e1, 'h1001a3, 'h1000e2, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h10003c, 'h2004f8, 'h100047, 'h1000e3, 'h1001b1, 'h1000e0, 'h1001b2, 'h1000e1, 'h1001b3, 'h1000e2, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h10003c, 'h2004f8, 'h100047, 'h1000e3, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1000e0, 'h1000e1, 'h1001c3, 'h1000e2, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h10003c, 'h2004f8, 'h100047, 'h1000e3, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000e0, 'h1000e1, 'h1001d3, 'h1000e2, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h10003c, 'h2004f8, 'h100047, 'h1000e3, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000e0, 'h1001e3, 'h1000e1, 'h1001e4, 'h1000e2, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h10003c, 'h2004f8, 'h100047, 'h1001e9, 'h1000e3, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000e0, 'h1001f3, 'h1000e1, 'h1001f4, 'h1000e2, 'h1001f5, 'h1001f6, 'h10003c, 'h2004f8, 'h100047, 'h1001f7, 'h1001f8, 'h1001f9, 'h1000e3, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h1000e0, 'h100203, 'h1000e1, 'h100204, 'h1000e2, 'h10003c, 'h2004f8, 'h100047, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h1000e3, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000e0, 'h100213, 'h1000e1, 'h10003c, 'h2004f8, 'h100047, 'h100214, 'h1000e2, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h1000e3, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000e0, 'h10003c, 'h2004f8, 'h100047, 'h100223, 'h1000e1, 'h100224, 'h1000e2, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h1000e3, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h10003c, 'h2004f8, 'h100047, 'h100232, 'h1000e0, 'h100233, 'h1000e1, 'h100234, 'h1000e2, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h1000e3, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h10003c, 'h2004f8, 'h100047, 'h100240, 'h100241, 'h100242, 'h100243, 'h1000e0, 'h1000e1, 'h100244, 'h1000e2, 'h100245, 'h100246, 'h100247, 'h1000e3, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10003c, 'h2004f8, 'h100047, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h1000e0, 'h1000e1, 'h100254, 'h1000e2, 'h100255, 'h1000e3, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10003c, 'h2004f8, 'h100047, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h1000e0, 'h100264, 'h1000e1, 'h100265, 'h1000e2, 'h100266, 'h1000e3, 'h100267, 'h100268, 'h100269, 'h10003c, 'h2004f8, 'h100047, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000e7, 'h1000e4, 'h100172, 'h1000e5, 'h100173, 'h1000e6, 'h100174, 'h100175, 'h10003c, 'h2004f8, 'h100047, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000e7, 'h100181, 'h1000e4, 'h100182, 'h1000e5, 'h100183, 'h1000e6, 'h10003c, 'h2004f8, 'h100047, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h100190, 'h1000e7, 'h100191, 'h1000e4, 'h100192, 'h1000e5, 'h10003c, 'h2004f8, 'h100047, 'h100193, 'h1000e6, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1000e7, 'h1001a1, 'h1000e4, 'h10003c, 'h2004f8, 'h100047, 'h1001a2, 'h1000e5, 'h1001a3, 'h1000e6, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1000e7, 'h10003c, 'h2004f8, 'h100047, 'h1001b1, 'h1001b2, 'h1000e4, 'h1000e5, 'h1001b3, 'h1000e6, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1000e7, 'h10003c, 'h2004f8, 'h100047, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1000e4, 'h1000e5, 'h1001c3, 'h1000e6, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1000e7, 'h10003c, 'h2004f8, 'h100047, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000e4, 'h1000e5, 'h1001d3, 'h1000e6, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1000e7, 'h10003c, 'h2004f8, 'h100047, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000e4, 'h1000e5, 'h1001e3, 'h1000e6, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1000e7, 'h10003c, 'h2004f8, 'h100047, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000e4, 'h1001f3, 'h1000e5, 'h1001f4, 'h1000e6, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h10003c, 'h2004f8, 'h100047, 'h1001f9, 'h1000e7, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h1000e4, 'h100203, 'h1000e5, 'h100204, 'h1000e6, 'h100205, 'h100206, 'h10003c, 'h2004f8, 'h100047, 'h100207, 'h100208, 'h100209, 'h1000e7, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000e4, 'h100213, 'h1000e5, 'h100214, 'h1000e6, 'h10003c, 'h2004f8, 'h100047, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h1000e7, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000e4, 'h100223, 'h1000e5, 'h10003c, 'h2004f8, 'h100047, 'h100224, 'h1000e6, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h1000e7, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h1000e4, 'h10003c, 'h2004f8, 'h100047, 'h1000e5, 'h100234, 'h1000e6, 'h100235, 'h100236, 'h100237, 'h1000e7, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h10003c, 'h2004f8, 'h100047, 'h100243, 'h1000e4, 'h1000e5, 'h100244, 'h1000e6, 'h100245, 'h1000e7, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h10003c, 'h2004f8, 'h100047, 'h100251, 'h100252, 'h100253, 'h1000e4, 'h1000e5, 'h100254, 'h1000e6, 'h100255, 'h1000e7, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10003c, 'h2004f8, 'h100047, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h1000e4, 'h1000e5, 'h100264, 'h1000e6, 'h100265, 'h1000e7, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10003c, 'h2004f8, 'h100047, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000eb, 'h1000e8, 'h100172, 'h1000e9, 'h100173, 'h1000ea, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h10003c, 'h2004f8, 'h100047, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000eb, 'h100181, 'h1000e8, 'h100182, 'h1000e9, 'h100183, 'h1000ea, 'h100184, 'h100185, 'h100186, 'h10003c, 'h2004f8, 'h100047, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h100190, 'h1000eb, 'h100191, 'h1000e8, 'h100192, 'h1000e9, 'h100193, 'h1000ea, 'h100194, 'h10003c, 'h2004f8, 'h100047, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1000eb, 'h1001a1, 'h1000e8, 'h1001a2, 'h1000e9, 'h1001a3, 'h10003c, 'h2004f8, 'h100047, 'h1000ea, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1000eb, 'h1001b1, 'h1001b2, 'h1000e8, 'h10003c, 'h2004f8, 'h100047, 'h1000e9, 'h1001b3, 'h1000ea, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1000eb, 'h1001bf, 'h1001c0, 'h1001c1, 'h10003c, 'h2004f8, 'h100047, 'h1001c2, 'h1000e8, 'h1000e9, 'h1001c3, 'h1000ea, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1000eb, 'h1001cd, 'h1001ce, 'h1001cf, 'h10003c, 'h2004f8, 'h100047, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000e8, 'h1000e9, 'h1001d3, 'h1000ea, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1000eb, 'h1001db, 'h1001dc, 'h1001dd, 'h10003c, 'h2004f8, 'h100047, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000e8, 'h1000e9, 'h1001e3, 'h1000ea, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1000eb, 'h1001e9, 'h1001ea, 'h1001eb, 'h10003c, 'h2004f8, 'h100047, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000e8, 'h1001f3, 'h1000e9, 'h1001f4, 'h1000ea, 'h1001f5, 'h1001f6, 'h1000eb, 'h1001f7, 'h1001f8, 'h1001f9, 'h10003c, 'h2004f8, 'h100047, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h1000e8, 'h100203, 'h1000e9, 'h100204, 'h1000ea, 'h100205, 'h1000eb, 'h100206, 'h100207, 'h10003c, 'h2004f8, 'h100047, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000e8, 'h100213, 'h1000e9, 'h100214, 'h1000ea, 'h100215, 'h1000eb, 'h10003c, 'h2004f8, 'h100047, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000e8, 'h100223, 'h1000e9, 'h100224, 'h1000ea, 'h10003c, 'h2004f8, 'h100047, 'h100225, 'h1000eb, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h1000e8, 'h1000e9, 'h10003c, 'h2004f8, 'h100047, 'h100234, 'h1000ea, 'h100235, 'h1000eb, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h10003c, 'h2004f8, 'h100047, 'h1000e8, 'h1000e9, 'h100244, 'h1000ea, 'h100245, 'h1000eb, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h10003c, 'h2004f8, 'h100047, 'h100252, 'h100253, 'h1000e8, 'h1000e9, 'h100254, 'h1000ea, 'h100255, 'h1000eb, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h10003c, 'h2004f8, 'h100047, 'h100260, 'h100261, 'h100262, 'h100263, 'h1000e8, 'h1000e9, 'h100264, 'h1000ea, 'h100265, 'h1000eb, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10003c, 'h2004f8, 'h100047, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000ef, 'h1000ec, 'h100172, 'h1000ed, 'h100173, 'h1000ee, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10003c, 'h2004f8, 'h100047, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000ef, 'h100181, 'h1000ec, 'h100182, 'h1000ed, 'h100183, 'h1000ee, 'h100184, 'h100185, 'h100186, 'h100187, 'h10003c, 'h2004f8, 'h100047, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h100190, 'h1000ef, 'h100191, 'h1000ec, 'h100192, 'h1000ed, 'h100193, 'h1000ee, 'h100194, 'h100195, 'h10003c, 'h2004f8, 'h100047, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1000ef, 'h1001a1, 'h1000ec, 'h1001a2, 'h1000ed, 'h1001a3, 'h1000ee, 'h10003c, 'h2004f8, 'h100047, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h1000ef, 'h1001b1, 'h1001b2, 'h1000ec, 'h1000ed, 'h1001b3, 'h10003c, 'h2004f8, 'h100047, 'h1000ee, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1000ef, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1000ec, 'h10003c, 'h2004f8, 'h100047, 'h1000ed, 'h1001c3, 'h1000ee, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1000ef, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h10003c, 'h2004f8, 'h100047, 'h1001d2, 'h1000ec, 'h1000ed, 'h1001d3, 'h1000ee, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1000ef, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h10003c, 'h2004f8, 'h100047, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000ec, 'h1000ed, 'h1001e3, 'h1000ee, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1000ef, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h10003c, 'h2004f8, 'h100047, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1000ec, 'h1001f3, 'h1000ed, 'h1001f4, 'h1000ee, 'h1001f5, 'h1001f6, 'h1000ef, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h10003c, 'h2004f8, 'h100047, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h1000ec, 'h100203, 'h1000ed, 'h100204, 'h1000ee, 'h100205, 'h1000ef, 'h100206, 'h100207, 'h100208, 'h100209, 'h10003c, 'h2004f8, 'h100047, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000ec, 'h100213, 'h1000ed, 'h100214, 'h1000ee, 'h100215, 'h1000ef, 'h100216, 'h100217, 'h10003c, 'h2004f8, 'h100047, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000ec, 'h100223, 'h1000ed, 'h100224, 'h1000ee, 'h100225, 'h1000ef, 'h10003c, 'h2004f8, 'h100047, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h1000ec, 'h1000ed, 'h100234, 'h1000ee, 'h100235, 'h10003c, 'h2004f8, 'h100047, 'h1000ef, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h1000ec, 'h1000ed, 'h100244, 'h10003c, 'h2004f8, 'h100047, 'h1000ee, 'h100245, 'h1000ef, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h1000ec, 'h10003c, 'h2004f8, 'h100047, 'h1000ed, 'h100254, 'h1000ee, 'h100255, 'h1000ef, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h10003c, 'h2004f8, 'h100047, 'h100263, 'h1000ec, 'h1000ed, 'h100264, 'h1000ee, 'h100265, 'h1000ef, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h10003c, 'h2004f8, 'h100047, 'h100271, 'h100272, 'h100171, 'h1000f3, 'h1000f0, 'h100172, 'h1000f1, 'h100173, 'h1000f2, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10003c, 'h2004f8, 'h100047, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000f3, 'h100181, 'h1000f0, 'h100182, 'h1000f1, 'h100183, 'h1000f2, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10003c, 'h2004f8, 'h100047, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h100190, 'h1000f3, 'h100191, 'h1000f0, 'h100192, 'h1000f1, 'h100193, 'h1000f2, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h10003c, 'h2004f8, 'h100047, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1000f3, 'h1001a1, 'h1000f0, 'h1001a2, 'h1000f1, 'h1001a3, 'h1000f2, 'h1001a4, 'h1001a5, 'h1001a6, 'h10003c, 'h2004f8, 'h100047, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h1000f3, 'h1001b1, 'h1001b2, 'h1000f0, 'h1000f1, 'h1001b3, 'h1000f2, 'h1001b4, 'h1001b5, 'h1001b6, 'h10003c, 'h2004f8, 'h100047, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1000f3, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1000f0, 'h1000f1, 'h1001c3, 'h1000f2, 'h1001c4, 'h10003c, 'h2004f8, 'h100047, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1000f3, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1000f0, 'h1000f1, 'h1001d3, 'h10003c, 'h2004f8, 'h100047, 'h1000f2, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1000f3, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1000f0, 'h10003c, 'h2004f8, 'h100047, 'h1000f1, 'h1001e3, 'h1000f2, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1000f3, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h10003c, 'h2004f8, 'h100047, 'h1001f2, 'h1000f0, 'h1001f3, 'h1000f1, 'h1001f4, 'h1000f2, 'h1001f5, 'h1001f6, 'h1000f3, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h10003c, 'h2004f8, 'h100047, 'h100200, 'h100201, 'h100202, 'h1000f0, 'h100203, 'h1000f1, 'h100204, 'h1000f2, 'h100205, 'h1000f3, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10003c, 'h2004f8, 'h100047, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h1000f0, 'h100213, 'h1000f1, 'h100214, 'h1000f2, 'h100215, 'h1000f3, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10003c, 'h2004f8, 'h100047, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h1000f0, 'h100223, 'h1000f1, 'h100224, 'h1000f2, 'h100225, 'h1000f3, 'h100226, 'h100227, 'h100228, 'h100229, 'h10003c, 'h2004f8, 'h100047, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h1000f0, 'h1000f1, 'h100234, 'h1000f2, 'h100235, 'h1000f3, 'h100236, 'h100237, 'h100238, 'h100239, 'h10003c, 'h2004f8, 'h100047, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h1000f0, 'h1000f1, 'h100244, 'h1000f2, 'h100245, 'h1000f3, 'h100246, 'h100247, 'h10003c, 'h2004f8, 'h100047, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h1000f0, 'h1000f1, 'h100254, 'h1000f2, 'h100255, 'h1000f3, 'h10003c, 'h2004f8, 'h100047, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f};
	int DATA3 [3*SIZE-1:0] = {DATA2, DATA0};
	
endpackage
