

package MATRIX_MULTIPLY_32_PKG_4;
	
	import MATRIX_MULTIPLY_32_PKG_3::DATA3;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h21f8d, 'h10803, 'h10957, 'h10813, 'h10823, 'h10958, 'h10833, 'h10843, 'h10959, 'h10b53, 'h10853, 'h10863, 'h1095a, 'h10873, 'h10883, 'h1095b, 'h103bc, 'h10893, 'h108a3, 'h1095c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b3, 'h108c3, 'h1095d, 'h108d3, 'h106e3, 'h1095e, 'h10b63, 'h106f3, 'h10703, 'h1095f, 'h10713, 'h10723, 'h10960, 'h10733, 'h103bc, 'h10743, 'h10961, 'h10753, 'h21f8e, 'h21f8f, 'h21f8d, 'h10763, 'h10962, 'h10773, 'h10783, 'h10963, 'h10793, 'h10b63, 'h107a3, 'h10964, 'h107b3, 'h107c3, 'h10965, 'h107d3, 'h107e3, 'h10966, 'h103bc, 'h107f3, 'h10803, 'h10967, 'h21f8e, 'h21f8f, 'h21f8d, 'h10813, 'h10823, 'h10968, 'h10833, 'h10843, 'h10969, 'h10b63, 'h10853, 'h10863, 'h1096a, 'h10873, 'h10883, 'h1096b, 'h10893, 'h103bc, 'h108a3, 'h1096c, 'h108b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c3, 'h1096d, 'h108d3, 'h106e3, 'h1096e, 'h10b73, 'h106f3, 'h10703, 'h1096f, 'h10713, 'h10723, 'h10970, 'h10733, 'h10743, 'h10971, 'h103bc, 'h10753, 'h10763, 'h10972, 'h21f8e, 'h21f8f, 'h21f8d, 'h10773, 'h10783, 'h10973, 'h10793, 'h10b73, 'h107a3, 'h10974, 'h107b3, 'h107c3, 'h10975, 'h107d3, 'h107e3, 'h10976, 'h107f3, 'h103bc, 'h10803, 'h10977, 'h10813, 'h21f8e, 'h21f8f, 'h21f8d, 'h10823, 'h10978, 'h10833, 'h10843, 'h10979, 'h10b73, 'h10853, 'h10863, 'h1097a, 'h10873, 'h10883, 'h1097b, 'h10893, 'h108a3, 'h1097c, 'h103bc, 'h108b3, 'h108c3, 'h1097d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d3, 'h106e3, 'h1097e, 'h10b83, 'h106f3, 'h10703, 'h1097f, 'h10713, 'h10723, 'h10980, 'h10733, 'h10743, 'h10981, 'h10753, 'h103bc, 'h10763, 'h10982, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10783, 'h10983, 'h10793, 'h10b83, 'h107a3, 'h10984, 'h107b3, 'h107c3, 'h10985, 'h107d3, 'h107e3, 'h10986, 'h107f3, 'h10803, 'h10987, 'h103bc, 'h10813, 'h10823, 'h10988, 'h21f8e, 'h21f8f, 'h21f8d, 'h10833, 'h10843, 'h10989, 'h10b83, 'h10853, 'h10863, 'h1098a, 'h10873, 'h10883, 'h1098b, 'h10893, 'h108a3, 'h1098c, 'h108b3, 'h103bc, 'h108c3, 'h1098d, 'h108d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1098e, 'h10b93, 'h106f3, 'h10703, 'h1098f, 'h10713, 'h10723, 'h10990, 'h10733, 'h10743, 'h10991, 'h10753, 'h10763, 'h10992, 'h103bc, 'h10773, 'h10783, 'h10993, 'h21f8e, 'h21f8f, 'h21f8d, 'h10793, 'h10b93, 'h107a3, 'h10994, 'h107b3, 'h107c3, 'h10995, 'h107d3, 'h107e3, 'h10996, 'h107f3, 'h10803, 'h10997, 'h10813, 'h103bc, 'h10823, 'h10998, 'h10833, 'h21f8e, 'h21f8f, 'h21f8d, 'h10843, 'h10999, 'h10b93, 'h10853, 'h10863, 'h1099a, 'h10873, 'h10883, 'h1099b, 'h10893, 'h108a3, 'h1099c, 'h108b3, 'h108c3, 'h1099d, 'h103bc, 'h108d3, 'h106e3, 'h1099e, 'h10ba3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f3, 'h10703, 'h1099f, 'h10713, 'h10723, 'h109a0, 'h10733, 'h10743, 'h109a1, 'h10753, 'h10763, 'h109a2, 'h10773, 'h103bc, 'h10783, 'h109a3, 'h10793, 'h10ba3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a3, 'h109a4, 'h107b3, 'h107c3, 'h109a5, 'h107d3, 'h107e3, 'h109a6, 'h107f3, 'h10803, 'h109a7, 'h10813, 'h10823, 'h109a8, 'h103bc, 'h10833, 'h10843, 'h109a9, 'h10ba3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10853, 'h10863, 'h109aa, 'h10873, 'h10883, 'h109ab, 'h10893, 'h108a3, 'h109ac, 'h108b3, 'h108c3, 'h109ad, 'h108d3, 'h103bc, 'h106e3, 'h109ae, 'h10bb3, 'h106f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10703, 'h109af, 'h10713, 'h10723, 'h109b0, 'h10733, 'h10743, 'h109b1, 'h10753, 'h10763, 'h109b2, 'h10773, 'h10783, 'h109b3, 'h103bc, 'h10793, 'h10bb3, 'h107a3, 'h109b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b3, 'h107c3, 'h109b5, 'h107d3, 'h107e3, 'h109b6, 'h107f3, 'h10803, 'h109b7, 'h10813, 'h10823, 'h109b8, 'h10833, 'h103bc, 'h10843, 'h109b9, 'h10bb3, 'h10853, 'h21f8e, 'h21f8f, 'h21f8d, 'h10863, 'h109ba, 'h10873, 'h10883, 'h109bb, 'h10893, 'h108a3, 'h109bc, 'h108b3, 'h108c3, 'h109bd, 'h108d3, 'h106e3, 'h109be, 'h10bc3, 'h103bc, 'h106f3, 'h10703, 'h109bf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10713, 'h10723, 'h109c0, 'h10733, 'h10743, 'h109c1, 'h10753, 'h10763, 'h109c2, 'h10773, 'h10783, 'h109c3, 'h10793, 'h10bc3, 'h103bc, 'h107a3, 'h109c4, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c3, 'h109c5, 'h107d3, 'h107e3, 'h109c6, 'h107f3, 'h10803, 'h109c7, 'h10813, 'h10823, 'h109c8, 'h10833, 'h10843, 'h109c9, 'h10bc3, 'h103bc, 'h10853, 'h10863, 'h109ca, 'h21f8e, 'h21f8f, 'h21f8d, 'h10873, 'h10883, 'h109cb, 'h10893, 'h108a3, 'h109cc, 'h108b3, 'h108c3, 'h109cd, 'h108d3, 'h106e3, 'h109ce, 'h10bd3, 'h106f3, 'h103bc, 'h10703, 'h109cf, 'h10713, 'h21f8e, 'h21f8f, 'h21f8d, 'h10723, 'h109d0, 'h10733, 'h10743, 'h109d1, 'h10753, 'h10763, 'h109d2, 'h10773, 'h10783, 'h109d3, 'h10793, 'h10bd3, 'h107a3, 'h109d4, 'h103bc, 'h107b3, 'h107c3, 'h109d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d3, 'h107e3, 'h109d6, 'h107f3, 'h10803, 'h109d7, 'h10813, 'h10823, 'h109d8, 'h10833, 'h10843, 'h109d9, 'h10bd3, 'h10853, 'h103bc, 'h10863, 'h109da, 'h10873, 'h21f8e, 'h21f8f, 'h21f8d, 'h10883, 'h109db, 'h10893, 'h108a3, 'h109dc, 'h108b3, 'h108c3, 'h109dd, 'h108d3, 'h106e3, 'h109de, 'h10be3, 'h106f3, 'h10703, 'h109df, 'h103bc, 'h10713, 'h10723, 'h109e0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10733, 'h10743, 'h109e1, 'h10753, 'h10763, 'h109e2, 'h10773, 'h10783, 'h109e3, 'h10793, 'h10be3, 'h107a3, 'h109e4, 'h107b3, 'h103bc, 'h107c3, 'h109e5, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e3, 'h109e6, 'h107f3, 'h10803, 'h109e7, 'h10813, 'h10823, 'h109e8, 'h10833, 'h10843, 'h109e9, 'h10be3, 'h10853, 'h10863, 'h109ea, 'h103bc, 'h10873, 'h10883, 'h109eb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10893, 'h108a3, 'h109ec, 'h108b3, 'h108c3, 'h109ed, 'h108d3, 'h106e3, 'h109ee, 'h10bf3, 'h106f3, 'h10703, 'h109ef, 'h10713, 'h103bc, 'h10723, 'h109f0, 'h10733, 'h21f8e, 'h21f8f, 'h21f8d, 'h10743, 'h109f1, 'h10753, 'h10763, 'h109f2, 'h10773, 'h10783, 'h109f3, 'h10793, 'h10bf3, 'h107a3, 'h109f4, 'h107b3, 'h107c3, 'h109f5, 'h103bc, 'h107d3, 'h107e3, 'h109f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f3, 'h10803, 'h109f7, 'h10813, 'h10823, 'h109f8, 'h10833, 'h10843, 'h109f9, 'h10bf3, 'h10853, 'h10863, 'h109fa, 'h10873, 'h103bc, 'h10883, 'h109fb, 'h10893, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a3, 'h109fc, 'h108b3, 'h108c3, 'h109fd, 'h108d3, 'h106e3, 'h109fe, 'h10c03, 'h106f3, 'h10703, 'h109ff, 'h10713, 'h10723, 'h10a00, 'h103bc, 'h10733, 'h10743, 'h10a01, 'h21f8e, 'h21f8f, 'h21f8d, 'h10753, 'h10763, 'h10a02, 'h10773, 'h10783, 'h10a03, 'h10793, 'h10c03, 'h107a3, 'h10a04, 'h107b3, 'h107c3, 'h10a05, 'h107d3, 'h103bc, 'h107e3, 'h10a06, 'h107f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10803, 'h10a07, 'h10813, 'h10823, 'h10a08, 'h10833, 'h10843, 'h10a09, 'h10c03, 'h10853, 'h10863, 'h10a0a, 'h10873, 'h10883, 'h10a0b, 'h103bc, 'h10893, 'h108a3, 'h10a0c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b3, 'h108c3, 'h10a0d, 'h108d3, 'h106e3, 'h10a0e, 'h10c13, 'h106f3, 'h10703, 'h10a0f, 'h10713, 'h10723, 'h10a10, 'h10733, 'h103bc, 'h10743, 'h10a11, 'h10753, 'h21f8e, 'h21f8f, 'h21f8d, 'h10763, 'h10a12, 'h10773, 'h10783, 'h10a13, 'h10793, 'h10c13, 'h107a3, 'h10a14, 'h107b3, 'h107c3, 'h10a15, 'h107d3, 'h107e3, 'h10a16, 'h103bc, 'h107f3, 'h10803, 'h10a17, 'h21f8e, 'h21f8f, 'h21f8d, 'h10813, 'h10823, 'h10a18, 'h10833, 'h10843, 'h10a19, 'h10c13, 'h10853, 'h10863, 'h10a1a, 'h10873, 'h10883, 'h10a1b, 'h10893, 'h103bc, 'h108a3, 'h10a1c, 'h108b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c3, 'h10a1d, 'h108d3, 'h106e3, 'h10a1e, 'h10c23, 'h106f3, 'h10703, 'h10a1f, 'h10713, 'h10723, 'h10a20, 'h10733, 'h10743, 'h10a21, 'h103bc, 'h10753, 'h10763, 'h10a22, 'h21f8e, 'h21f8f, 'h21f8d, 'h10773, 'h10783, 'h10a23, 'h10793, 'h10c23, 'h107a3, 'h10a24, 'h107b3, 'h107c3, 'h10a25, 'h107d3, 'h107e3, 'h10a26, 'h107f3, 'h103bc, 'h10803, 'h10a27, 'h10813, 'h21f8e, 'h21f8f, 'h21f8d, 'h10823, 'h10a28, 'h10833, 'h10843, 'h10a29, 'h10c23, 'h10853, 'h10863, 'h10a2a, 'h10873, 'h10883, 'h10a2b, 'h10893, 'h108a3, 'h10a2c, 'h103bc, 'h108b3, 'h108c3, 'h10a2d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d3, 'h106e3, 'h10a2e, 'h10c33, 'h106f3, 'h10703, 'h10a2f, 'h10713, 'h10723, 'h10a30, 'h10733, 'h10743, 'h10a31, 'h10753, 'h103bc, 'h10763, 'h10a32, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10783, 'h10a33, 'h10793, 'h10c33, 'h107a3, 'h10a34, 'h107b3, 'h107c3, 'h10a35, 'h107d3, 'h107e3, 'h10a36, 'h107f3, 'h10803, 'h10a37, 'h103bc, 'h10813, 'h10823, 'h10a38, 'h21f8e, 'h21f8f, 'h21f8d, 'h10833, 'h10843, 'h10a39, 'h10c33, 'h10853, 'h10863, 'h10a3a, 'h10873, 'h10883, 'h10a3b, 'h10893, 'h108a3, 'h10a3c, 'h108b3, 'h103bc, 'h108c3, 'h10a3d, 'h108d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h10a3e, 'h10c43, 'h106f3, 'h10703, 'h10a3f, 'h10713, 'h10723, 'h10a40, 'h10733, 'h10743, 'h10a41, 'h10753, 'h10763, 'h10a42, 'h103bc, 'h10773, 'h10783, 'h10a43, 'h21f8e, 'h21f8f, 'h21f8d, 'h10793, 'h10c43, 'h107a3, 'h10a44, 'h107b3, 'h107c3, 'h10a45, 'h107d3, 'h107e3, 'h10a46, 'h107f3, 'h10803, 'h10a47, 'h10813, 'h103bc, 'h10823, 'h10a48, 'h10833, 'h21f8e, 'h21f8f, 'h21f8d, 'h10843, 'h10a49, 'h10c43, 'h10853, 'h10863, 'h10a4a, 'h10873, 'h10883, 'h10a4b, 'h10893, 'h108a3, 'h10a4c, 'h108b3, 'h108c3, 'h10a4d, 'h103bc, 'h108d3, 'h106e3, 'h10a4e, 'h10c53, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f3, 'h10703, 'h10a4f, 'h10713, 'h10723, 'h10a50, 'h10733, 'h10743, 'h10a51, 'h10753, 'h10763, 'h10a52, 'h10773, 'h103bc, 'h10783, 'h10a53, 'h10793, 'h10c53, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a3, 'h10a54, 'h107b3, 'h107c3, 'h10a55, 'h107d3, 'h107e3, 'h10a56, 'h107f3, 'h10803, 'h10a57, 'h10813, 'h10823, 'h10a58, 'h103bc, 'h10833, 'h10843, 'h10a59, 'h10c53, 'h21f8e, 'h21f8f, 'h21f8d, 'h10853, 'h10863, 'h10a5a, 'h10873, 'h10883, 'h10a5b, 'h10893, 'h108a3, 'h10a5c, 'h108b3, 'h108c3, 'h10a5d, 'h108d3, 'h103bc, 'h106e3, 'h10a5e, 'h10c63, 'h106f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10703, 'h10a5f, 'h10713, 'h10723, 'h10a60, 'h10733, 'h10743, 'h10a61, 'h10753, 'h10763, 'h10a62, 'h10773, 'h10783, 'h10a63, 'h103bc, 'h10793, 'h10c63, 'h107a3, 'h10a64, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b3, 'h107c3, 'h10a65, 'h107d3, 'h107e3, 'h10a66, 'h107f3, 'h10803, 'h10a67, 'h10813, 'h10823, 'h10a68, 'h10833, 'h103bc, 'h10843, 'h10a69, 'h10c63, 'h10853, 'h21f8e, 'h21f8f, 'h21f8d, 'h10863, 'h10a6a, 'h10873, 'h10883, 'h10a6b, 'h10893, 'h108a3, 'h10a6c, 'h108b3, 'h108c3, 'h10a6d, 'h108d3, 'h106e3, 'h10a6e, 'h10c73, 'h103bc, 'h106f3, 'h10703, 'h10a6f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10713, 'h10723, 'h10a70, 'h10733, 'h10743, 'h10a71, 'h10753, 'h10763, 'h10a72, 'h10773, 'h10783, 'h10a73, 'h10793, 'h10c73, 'h103bc, 'h107a3, 'h10a74, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c3, 'h10a75, 'h107d3, 'h107e3, 'h10a76, 'h107f3, 'h10803, 'h10a77, 'h10813, 'h10823, 'h10a78, 'h10833, 'h10843, 'h10a79, 'h10c73, 'h103bc, 'h10853, 'h10863, 'h10a7a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10873, 'h10883, 'h10a7b, 'h10893, 'h108a3, 'h10a7c, 'h108b3, 'h108c3, 'h10a7d, 'h108d3, 'h106e3, 'h10a7e, 'h10c83, 'h106f3, 'h103bc, 'h10703, 'h10a7f, 'h10713, 'h21f8e, 'h21f8f, 'h21f8d, 'h10723, 'h10a80, 'h10733, 'h10743, 'h10a81, 'h10753, 'h10763, 'h10a82, 'h10773, 'h10783, 'h10a83, 'h10793, 'h10c83, 'h107a3, 'h10a84, 'h103bc, 'h107b3, 'h107c3, 'h10a85, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d3, 'h107e3, 'h10a86, 'h107f3, 'h10803, 'h10a87, 'h10813, 'h10823, 'h10a88, 'h10833, 'h10843, 'h10a89, 'h10c83, 'h10853, 'h103bc, 'h10863, 'h10a8a, 'h10873, 'h21f8e, 'h21f8f, 'h21f8d, 'h10883, 'h10a8b, 'h10893, 'h108a3, 'h10a8c, 'h108b3, 'h108c3, 'h10a8d, 'h108d3, 'h106e3, 'h10a8e, 'h10c93, 'h106f3, 'h10703, 'h10a8f, 'h103bc, 'h10713, 'h10723, 'h10a90, 'h21f8e, 'h21f8f, 'h21f8d, 'h10733, 'h10743, 'h10a91, 'h10753, 'h10763, 'h10a92, 'h10773, 'h10783, 'h10a93, 'h10793, 'h10c93, 'h107a3, 'h10a94, 'h107b3, 'h103bc, 'h107c3, 'h10a95, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e3, 'h10a96, 'h107f3, 'h10803, 'h10a97, 'h10813, 'h10823, 'h10a98, 'h10833, 'h10843, 'h10a99, 'h10c93, 'h10853, 'h10863, 'h10a9a, 'h103bc, 'h10873, 'h10883, 'h10a9b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10893, 'h108a3, 'h10a9c, 'h108b3, 'h108c3, 'h10a9d, 'h108d3, 'h106e3, 'h10a9e, 'h10ca3, 'h106f3, 'h10703, 'h10a9f, 'h10713, 'h103bc, 'h10723, 'h10aa0, 'h10733, 'h21f8e, 'h21f8f, 'h21f8d, 'h10743, 'h10aa1, 'h10753, 'h10763, 'h10aa2, 'h10773, 'h10783, 'h10aa3, 'h10793, 'h10ca3, 'h107a3, 'h10aa4, 'h107b3, 'h107c3, 'h10aa5, 'h103bc, 'h107d3, 'h107e3, 'h10aa6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f3, 'h10803, 'h10aa7, 'h10813, 'h10823, 'h10aa8, 'h10833, 'h10843, 'h10aa9, 'h10ca3, 'h10853, 'h10863, 'h10aaa, 'h10873, 'h103bc, 'h10883, 'h10aab, 'h10893, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a3, 'h10aac, 'h108b3, 'h108c3, 'h10aad, 'h108d3, 'h106e3, 'h10aae, 'h10cb3, 'h106f3, 'h10703, 'h10aaf, 'h10713, 'h10723, 'h10ab0, 'h103bc, 'h10733, 'h10743, 'h10ab1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10753, 'h10763, 'h10ab2, 'h10773, 'h10783, 'h10ab3, 'h10793, 'h10cb3, 'h107a3, 'h10ab4, 'h107b3, 'h107c3, 'h10ab5, 'h107d3, 'h103bc, 'h107e3, 'h10ab6, 'h107f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10803, 'h10ab7, 'h10813, 'h10823, 'h10ab8, 'h10833, 'h10843, 'h10ab9, 'h10cb3, 'h10853, 'h10863, 'h10aba, 'h10873, 'h10883, 'h10abb, 'h103bc, 'h10893, 'h108a3, 'h10abc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b3, 'h108c3, 'h10abd, 'h108d3, 'h106e3, 'h10abe, 'h10cc3, 'h106f3, 'h10703, 'h10abf, 'h10713, 'h10723, 'h10ac0, 'h10733, 'h103bc, 'h10743, 'h10ac1, 'h10753, 'h21f8e, 'h21f8f, 'h21f8d, 'h10763, 'h10ac2, 'h10773, 'h10783, 'h10ac3, 'h10793, 'h10cc3, 'h107a3, 'h10ac4, 'h107b3, 'h107c3, 'h10ac5, 'h107d3, 'h107e3, 'h10ac6, 'h103bc, 'h107f3, 'h10803, 'h10ac7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10813, 'h10823, 'h10ac8, 'h10833, 'h10843, 'h10ac9, 'h10cc3, 'h10853, 'h10863, 'h10aca, 'h10873, 'h10883, 'h10acb, 'h10893, 'h103bc, 'h108a3, 'h10acc, 'h108b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c3, 'h10acd, 'h108d3, 'h106e3, 'h10ace, 'h10cd3, 'h106f3, 'h10703, 'h10acf, 'h10713, 'h10723, 'h10ad0, 'h10733, 'h10743, 'h10ad1, 'h103bc, 'h10753, 'h10763, 'h10ad2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10773, 'h10783, 'h10ad3, 'h10793, 'h10cd3, 'h107a3, 'h10ad4, 'h107b3, 'h107c3, 'h10ad5, 'h107d3, 'h107e3, 'h10ad6, 'h107f3, 'h103bc, 'h10803, 'h10ad7, 'h10813, 'h21f8e, 'h21f8f, 'h21f8d, 'h10823, 'h10ad8, 'h10833, 'h10843, 'h10ad9, 'h10cd3, 'h10853, 'h10863, 'h10ada, 'h10873, 'h10883, 'h10adb, 'h10893, 'h108a3, 'h10adc, 'h103bc, 'h108b3, 'h108c3, 'h10add, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d3, 'h106e4, 'h108de, 'h10ae4, 'h106f4, 'h10704, 'h108df, 'h10714, 'h10724, 'h108e0, 'h10734, 'h10744, 'h108e1, 'h10754, 'h103bc, 'h10764, 'h108e2, 'h10774, 'h21f8e, 'h21f8f, 'h21f8d, 'h10784, 'h108e3, 'h10794, 'h10ae4, 'h107a4, 'h108e4, 'h107b4, 'h107c4, 'h108e5, 'h107d4, 'h107e4, 'h108e6, 'h107f4, 'h10804, 'h108e7, 'h103bc, 'h10814, 'h10824, 'h108e8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10834, 'h10844, 'h108e9, 'h10ae4, 'h10854, 'h10864, 'h108ea, 'h10874, 'h10884, 'h108eb, 'h10894, 'h108a4, 'h108ec, 'h108b4, 'h103bc, 'h108c4, 'h108ed, 'h108d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h108ee, 'h10af4, 'h106f4, 'h10704, 'h108ef, 'h10714, 'h10724, 'h108f0, 'h10734, 'h10744, 'h108f1, 'h10754, 'h10764, 'h108f2, 'h103bc, 'h10774, 'h10784, 'h108f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10794, 'h10af4, 'h107a4, 'h108f4, 'h107b4, 'h107c4, 'h108f5, 'h107d4, 'h107e4, 'h108f6, 'h107f4, 'h10804, 'h108f7, 'h10814, 'h103bc, 'h10824, 'h108f8, 'h10834, 'h21f8e, 'h21f8f, 'h21f8d, 'h10844, 'h108f9, 'h10af4, 'h10854, 'h10864, 'h108fa, 'h10874, 'h10884, 'h108fb, 'h10894, 'h108a4, 'h108fc, 'h108b4, 'h108c4, 'h108fd, 'h103bc, 'h108d4, 'h106e4, 'h108fe, 'h10b04, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f4, 'h10704, 'h108ff, 'h10714, 'h10724, 'h10900, 'h10734, 'h10744, 'h10901, 'h10754, 'h10764, 'h10902, 'h10774, 'h103bc, 'h10784, 'h10903, 'h10794, 'h10b04, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a4, 'h10904, 'h107b4, 'h107c4, 'h10905, 'h107d4, 'h107e4, 'h10906, 'h107f4, 'h10804, 'h10907, 'h10814, 'h10824, 'h10908, 'h103bc, 'h10834, 'h10844, 'h10909, 'h10b04, 'h21f8e, 'h21f8f, 'h21f8d, 'h10854, 'h10864, 'h1090a, 'h10874, 'h10884, 'h1090b, 'h10894, 'h108a4, 'h1090c, 'h108b4, 'h108c4, 'h1090d, 'h108d4, 'h103bc, 'h106e4, 'h1090e, 'h10b14, 'h106f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10704, 'h1090f, 'h10714, 'h10724, 'h10910, 'h10734, 'h10744, 'h10911, 'h10754, 'h10764, 'h10912, 'h10774, 'h10784, 'h10913, 'h103bc, 'h10794, 'h10b14, 'h107a4, 'h10914, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b4, 'h107c4, 'h10915, 'h107d4, 'h107e4, 'h10916, 'h107f4, 'h10804, 'h10917, 'h10814, 'h10824, 'h10918, 'h10834, 'h103bc, 'h10844, 'h10919, 'h10b14, 'h10854, 'h21f8e, 'h21f8f, 'h21f8d, 'h10864, 'h1091a, 'h10874, 'h10884, 'h1091b, 'h10894, 'h108a4, 'h1091c, 'h108b4, 'h108c4, 'h1091d, 'h108d4, 'h106e4, 'h1091e, 'h10b24, 'h103bc, 'h106f4, 'h10704, 'h1091f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10714, 'h10724, 'h10920, 'h10734, 'h10744, 'h10921, 'h10754, 'h10764, 'h10922, 'h10774, 'h10784, 'h10923, 'h10794, 'h10b24, 'h103bc, 'h107a4, 'h10924, 'h107b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c4, 'h10925, 'h107d4, 'h107e4, 'h10926, 'h107f4, 'h10804, 'h10927, 'h10814, 'h10824, 'h10928, 'h10834, 'h10844, 'h10929, 'h10b24, 'h103bc, 'h10854, 'h10864, 'h1092a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10874, 'h10884, 'h1092b, 'h10894, 'h108a4, 'h1092c, 'h108b4, 'h108c4, 'h1092d, 'h108d4, 'h106e4, 'h1092e, 'h10b34, 'h106f4, 'h103bc, 'h10704, 'h1092f, 'h10714, 'h21f8e, 'h21f8f, 'h21f8d, 'h10724, 'h10930, 'h10734, 'h10744, 'h10931, 'h10754, 'h10764, 'h10932, 'h10774, 'h10784, 'h10933, 'h10794, 'h10b34, 'h107a4, 'h10934, 'h103bc, 'h107b4, 'h107c4, 'h10935, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d4, 'h107e4, 'h10936, 'h107f4, 'h10804, 'h10937, 'h10814, 'h10824, 'h10938, 'h10834, 'h10844, 'h10939, 'h10b34, 'h10854, 'h103bc, 'h10864, 'h1093a, 'h10874, 'h21f8e, 'h21f8f, 'h21f8d, 'h10884, 'h1093b, 'h10894, 'h108a4, 'h1093c, 'h108b4, 'h108c4, 'h1093d, 'h108d4, 'h106e4, 'h1093e, 'h10b44, 'h106f4, 'h10704, 'h1093f, 'h103bc, 'h10714, 'h10724, 'h10940, 'h21f8e, 'h21f8f, 'h21f8d, 'h10734, 'h10744, 'h10941, 'h10754, 'h10764, 'h10942, 'h10774, 'h10784, 'h10943, 'h10794, 'h10b44, 'h107a4, 'h10944, 'h107b4, 'h103bc, 'h107c4, 'h10945, 'h107d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e4, 'h10946, 'h107f4, 'h10804, 'h10947, 'h10814, 'h10824, 'h10948, 'h10834, 'h10844, 'h10949, 'h10b44, 'h10854, 'h10864, 'h1094a, 'h103bc, 'h10874, 'h10884, 'h1094b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10894, 'h108a4, 'h1094c, 'h108b4, 'h108c4, 'h1094d, 'h108d4, 'h106e4, 'h1094e, 'h10b54, 'h106f4, 'h10704, 'h1094f, 'h10714, 'h103bc, 'h10724, 'h10950, 'h10734, 'h21f8e, 'h21f8f, 'h21f8d, 'h10744, 'h10951, 'h10754, 'h10764, 'h10952, 'h10774, 'h10784, 'h10953, 'h10794, 'h10b54, 'h107a4, 'h10954, 'h107b4, 'h107c4, 'h10955, 'h103bc, 'h107d4, 'h107e4, 'h10956, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f4, 'h10804, 'h10957, 'h10814, 'h10824, 'h10958, 'h10834, 'h10844, 'h10959, 'h10b54, 'h10854, 'h10864, 'h1095a, 'h10874, 'h103bc, 'h10884, 'h1095b, 'h10894, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a4, 'h1095c, 'h108b4, 'h108c4, 'h1095d, 'h108d4, 'h106e4, 'h1095e, 'h10b64, 'h106f4, 'h10704, 'h1095f, 'h10714, 'h10724, 'h10960, 'h103bc, 'h10734, 'h10744, 'h10961, 'h21f8e, 'h21f8f, 'h21f8d, 'h10754, 'h10764, 'h10962, 'h10774, 'h10784, 'h10963, 'h10794, 'h10b64, 'h107a4, 'h10964, 'h107b4, 'h107c4, 'h10965, 'h107d4, 'h103bc, 'h107e4, 'h10966, 'h107f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10804, 'h10967, 'h10814, 'h10824, 'h10968, 'h10834, 'h10844, 'h10969, 'h10b64, 'h10854, 'h10864, 'h1096a, 'h10874, 'h10884, 'h1096b, 'h103bc, 'h10894, 'h108a4, 'h1096c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b4, 'h108c4, 'h1096d, 'h108d4, 'h106e4, 'h1096e, 'h10b74, 'h106f4, 'h10704, 'h1096f, 'h10714, 'h10724, 'h10970, 'h10734, 'h103bc, 'h10744, 'h10971, 'h10754, 'h21f8e, 'h21f8f, 'h21f8d, 'h10764, 'h10972, 'h10774, 'h10784, 'h10973, 'h10794, 'h10b74, 'h107a4, 'h10974, 'h107b4, 'h107c4, 'h10975, 'h107d4, 'h107e4, 'h10976, 'h103bc, 'h107f4, 'h10804, 'h10977, 'h21f8e, 'h21f8f, 'h21f8d, 'h10814, 'h10824, 'h10978, 'h10834, 'h10844, 'h10979, 'h10b74, 'h10854, 'h10864, 'h1097a, 'h10874, 'h10884, 'h1097b, 'h10894, 'h103bc, 'h108a4, 'h1097c, 'h108b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c4, 'h1097d, 'h108d4, 'h106e4, 'h1097e, 'h10b84, 'h106f4, 'h10704, 'h1097f, 'h10714, 'h10724, 'h10980, 'h10734, 'h10744, 'h10981, 'h103bc, 'h10754, 'h10764, 'h10982, 'h21f8e, 'h21f8f, 'h21f8d, 'h10774, 'h10784, 'h10983, 'h10794, 'h10b84, 'h107a4, 'h10984, 'h107b4, 'h107c4, 'h10985, 'h107d4, 'h107e4, 'h10986, 'h107f4, 'h103bc, 'h10804, 'h10987, 'h10814, 'h21f8e, 'h21f8f, 'h21f8d, 'h10824, 'h10988, 'h10834, 'h10844, 'h10989, 'h10b84, 'h10854, 'h10864, 'h1098a, 'h10874, 'h10884, 'h1098b, 'h10894, 'h108a4, 'h1098c, 'h103bc, 'h108b4, 'h108c4, 'h1098d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d4, 'h106e4, 'h1098e, 'h10b94, 'h106f4, 'h10704, 'h1098f, 'h10714, 'h10724, 'h10990, 'h10734, 'h10744, 'h10991, 'h10754, 'h103bc, 'h10764, 'h10992, 'h10774, 'h21f8e, 'h21f8f, 'h21f8d, 'h10784, 'h10993, 'h10794, 'h10b94, 'h107a4, 'h10994, 'h107b4, 'h107c4, 'h10995, 'h107d4, 'h107e4, 'h10996, 'h107f4, 'h10804, 'h10997, 'h103bc, 'h10814, 'h10824, 'h10998, 'h21f8e, 'h21f8f, 'h21f8d, 'h10834, 'h10844, 'h10999, 'h10b94, 'h10854, 'h10864, 'h1099a, 'h10874, 'h10884, 'h1099b, 'h10894, 'h108a4, 'h1099c, 'h108b4, 'h103bc, 'h108c4, 'h1099d, 'h108d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1099e, 'h10ba4, 'h106f4, 'h10704, 'h1099f, 'h10714, 'h10724, 'h109a0, 'h10734, 'h10744, 'h109a1, 'h10754, 'h10764, 'h109a2, 'h103bc, 'h10774, 'h10784, 'h109a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10794, 'h10ba4, 'h107a4, 'h109a4, 'h107b4, 'h107c4, 'h109a5, 'h107d4, 'h107e4, 'h109a6, 'h107f4, 'h10804, 'h109a7, 'h10814, 'h103bc, 'h10824, 'h109a8, 'h10834, 'h21f8e, 'h21f8f, 'h21f8d, 'h10844, 'h109a9, 'h10ba4, 'h10854, 'h10864, 'h109aa, 'h10874, 'h10884, 'h109ab, 'h10894, 'h108a4, 'h109ac, 'h108b4, 'h108c4, 'h109ad, 'h103bc, 'h108d4, 'h106e4, 'h109ae, 'h10bb4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f4, 'h10704, 'h109af, 'h10714, 'h10724, 'h109b0, 'h10734, 'h10744, 'h109b1, 'h10754, 'h10764, 'h109b2, 'h10774, 'h103bc, 'h10784, 'h109b3, 'h10794, 'h10bb4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a4, 'h109b4, 'h107b4, 'h107c4, 'h109b5, 'h107d4, 'h107e4, 'h109b6, 'h107f4, 'h10804, 'h109b7, 'h10814, 'h10824, 'h109b8, 'h103bc, 'h10834, 'h10844, 'h109b9, 'h10bb4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10854, 'h10864, 'h109ba, 'h10874, 'h10884, 'h109bb, 'h10894, 'h108a4, 'h109bc, 'h108b4, 'h108c4, 'h109bd, 'h108d4, 'h103bc, 'h106e4, 'h109be, 'h10bc4, 'h106f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10704, 'h109bf, 'h10714, 'h10724, 'h109c0, 'h10734, 'h10744, 'h109c1, 'h10754, 'h10764, 'h109c2, 'h10774, 'h10784, 'h109c3, 'h103bc, 'h10794, 'h10bc4, 'h107a4, 'h109c4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b4, 'h107c4, 'h109c5, 'h107d4, 'h107e4, 'h109c6, 'h107f4, 'h10804, 'h109c7, 'h10814, 'h10824, 'h109c8, 'h10834, 'h103bc, 'h10844, 'h109c9, 'h10bc4, 'h10854, 'h21f8e, 'h21f8f, 'h21f8d, 'h10864, 'h109ca, 'h10874, 'h10884, 'h109cb, 'h10894, 'h108a4, 'h109cc, 'h108b4, 'h108c4, 'h109cd, 'h108d4, 'h106e4, 'h109ce, 'h10bd4, 'h103bc, 'h106f4, 'h10704, 'h109cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10714, 'h10724, 'h109d0, 'h10734, 'h10744, 'h109d1, 'h10754, 'h10764, 'h109d2, 'h10774, 'h10784, 'h109d3, 'h10794, 'h10bd4, 'h103bc, 'h107a4, 'h109d4, 'h107b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c4, 'h109d5, 'h107d4, 'h107e4, 'h109d6, 'h107f4, 'h10804, 'h109d7, 'h10814, 'h10824, 'h109d8, 'h10834, 'h10844, 'h109d9, 'h10bd4, 'h103bc, 'h10854, 'h10864, 'h109da, 'h21f8e, 'h21f8f, 'h21f8d, 'h10874, 'h10884, 'h109db, 'h10894, 'h108a4, 'h109dc, 'h108b4, 'h108c4, 'h109dd, 'h108d4, 'h106e4, 'h109de, 'h10be4, 'h106f4, 'h103bc, 'h10704, 'h109df, 'h10714, 'h21f8e, 'h21f8f, 'h21f8d, 'h10724, 'h109e0, 'h10734, 'h10744, 'h109e1, 'h10754, 'h10764, 'h109e2, 'h10774, 'h10784, 'h109e3, 'h10794, 'h10be4, 'h107a4, 'h109e4, 'h103bc, 'h107b4, 'h107c4, 'h109e5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d4, 'h107e4, 'h109e6, 'h107f4, 'h10804, 'h109e7, 'h10814, 'h10824, 'h109e8, 'h10834, 'h10844, 'h109e9, 'h10be4, 'h10854, 'h103bc, 'h10864, 'h109ea, 'h10874, 'h21f8e, 'h21f8f, 'h21f8d, 'h10884, 'h109eb, 'h10894, 'h108a4, 'h109ec, 'h108b4, 'h108c4, 'h109ed, 'h108d4, 'h106e4, 'h109ee, 'h10bf4, 'h106f4, 'h10704, 'h109ef, 'h103bc, 'h10714, 'h10724, 'h109f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10734, 'h10744, 'h109f1, 'h10754, 'h10764, 'h109f2, 'h10774, 'h10784, 'h109f3, 'h10794, 'h10bf4, 'h107a4, 'h109f4, 'h107b4, 'h103bc, 'h107c4, 'h109f5, 'h107d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e4, 'h109f6, 'h107f4, 'h10804, 'h109f7, 'h10814, 'h10824, 'h109f8, 'h10834, 'h10844, 'h109f9, 'h10bf4, 'h10854, 'h10864, 'h109fa, 'h103bc, 'h10874, 'h10884, 'h109fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10894, 'h108a4, 'h109fc, 'h108b4, 'h108c4, 'h109fd, 'h108d4, 'h106e4, 'h109fe, 'h10c04, 'h106f4, 'h10704, 'h109ff, 'h10714, 'h103bc, 'h10724, 'h10a00, 'h10734, 'h21f8e, 'h21f8f, 'h21f8d, 'h10744, 'h10a01, 'h10754, 'h10764, 'h10a02, 'h10774, 'h10784, 'h10a03, 'h10794, 'h10c04, 'h107a4, 'h10a04, 'h107b4, 'h107c4, 'h10a05, 'h103bc, 'h107d4, 'h107e4, 'h10a06, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f4, 'h10804, 'h10a07, 'h10814, 'h10824, 'h10a08, 'h10834, 'h10844, 'h10a09, 'h10c04, 'h10854, 'h10864, 'h10a0a, 'h10874, 'h103bc, 'h10884, 'h10a0b, 'h10894, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a4, 'h10a0c, 'h108b4, 'h108c4, 'h10a0d, 'h108d4, 'h106e4, 'h10a0e, 'h10c14, 'h106f4, 'h10704, 'h10a0f, 'h10714, 'h10724, 'h10a10, 'h103bc, 'h10734, 'h10744, 'h10a11, 'h21f8e, 'h21f8f, 'h21f8d, 'h10754, 'h10764, 'h10a12, 'h10774, 'h10784, 'h10a13, 'h10794, 'h10c14, 'h107a4, 'h10a14, 'h107b4, 'h107c4, 'h10a15, 'h107d4, 'h103bc, 'h107e4, 'h10a16, 'h107f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10804, 'h10a17, 'h10814, 'h10824, 'h10a18, 'h10834, 'h10844, 'h10a19, 'h10c14, 'h10854, 'h10864, 'h10a1a, 'h10874, 'h10884, 'h10a1b, 'h103bc, 'h10894, 'h108a4, 'h10a1c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b4, 'h108c4, 'h10a1d, 'h108d4, 'h106e4, 'h10a1e, 'h10c24, 'h106f4, 'h10704, 'h10a1f, 'h10714, 'h10724, 'h10a20, 'h10734, 'h103bc, 'h10744, 'h10a21, 'h10754, 'h21f8e, 'h21f8f, 'h21f8d, 'h10764, 'h10a22, 'h10774, 'h10784, 'h10a23, 'h10794, 'h10c24, 'h107a4, 'h10a24, 'h107b4, 'h107c4, 'h10a25, 'h107d4, 'h107e4, 'h10a26, 'h103bc, 'h107f4, 'h10804, 'h10a27, 'h21f8e, 'h21f8f, 'h21f8d, 'h10814, 'h10824, 'h10a28, 'h10834, 'h10844, 'h10a29, 'h10c24, 'h10854, 'h10864, 'h10a2a, 'h10874, 'h10884, 'h10a2b, 'h10894, 'h103bc, 'h108a4, 'h10a2c, 'h108b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c4, 'h10a2d, 'h108d4, 'h106e4, 'h10a2e, 'h10c34, 'h106f4, 'h10704, 'h10a2f, 'h10714, 'h10724, 'h10a30, 'h10734, 'h10744, 'h10a31, 'h103bc, 'h10754, 'h10764, 'h10a32, 'h21f8e, 'h21f8f, 'h21f8d, 'h10774, 'h10784, 'h10a33, 'h10794, 'h10c34, 'h107a4, 'h10a34, 'h107b4, 'h107c4, 'h10a35, 'h107d4, 'h107e4, 'h10a36, 'h107f4, 'h103bc, 'h10804, 'h10a37, 'h10814, 'h21f8e, 'h21f8f, 'h21f8d, 'h10824, 'h10a38, 'h10834, 'h10844, 'h10a39, 'h10c34, 'h10854, 'h10864, 'h10a3a, 'h10874, 'h10884, 'h10a3b, 'h10894, 'h108a4, 'h10a3c, 'h103bc, 'h108b4, 'h108c4, 'h10a3d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d4, 'h106e4, 'h10a3e, 'h10c44, 'h106f4, 'h10704, 'h10a3f, 'h10714, 'h10724, 'h10a40, 'h10734, 'h10744, 'h10a41, 'h10754, 'h103bc, 'h10764, 'h10a42, 'h10774, 'h21f8e, 'h21f8f, 'h21f8d, 'h10784, 'h10a43, 'h10794, 'h10c44, 'h107a4, 'h10a44, 'h107b4, 'h107c4, 'h10a45, 'h107d4, 'h107e4, 'h10a46, 'h107f4, 'h10804, 'h10a47, 'h103bc, 'h10814, 'h10824, 'h10a48, 'h21f8e, 'h21f8f, 'h21f8d, 'h10834, 'h10844, 'h10a49, 'h10c44, 'h10854, 'h10864, 'h10a4a, 'h10874, 'h10884, 'h10a4b, 'h10894, 'h108a4, 'h10a4c, 'h108b4, 'h103bc, 'h108c4, 'h10a4d, 'h108d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h10a4e, 'h10c54, 'h106f4, 'h10704, 'h10a4f, 'h10714, 'h10724, 'h10a50, 'h10734, 'h10744, 'h10a51, 'h10754, 'h10764, 'h10a52, 'h103bc, 'h10774, 'h10784, 'h10a53, 'h21f8e, 'h21f8f, 'h21f8d, 'h10794, 'h10c54, 'h107a4, 'h10a54, 'h107b4, 'h107c4, 'h10a55, 'h107d4, 'h107e4, 'h10a56, 'h107f4, 'h10804, 'h10a57, 'h10814, 'h103bc, 'h10824, 'h10a58, 'h10834, 'h21f8e, 'h21f8f, 'h21f8d, 'h10844, 'h10a59, 'h10c54, 'h10854, 'h10864, 'h10a5a, 'h10874, 'h10884, 'h10a5b, 'h10894, 'h108a4, 'h10a5c, 'h108b4, 'h108c4, 'h10a5d, 'h103bc, 'h108d4, 'h106e4, 'h10a5e, 'h10c64, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f4, 'h10704, 'h10a5f, 'h10714, 'h10724, 'h10a60, 'h10734, 'h10744, 'h10a61, 'h10754, 'h10764, 'h10a62, 'h10774, 'h103bc, 'h10784, 'h10a63, 'h10794, 'h10c64, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a4, 'h10a64, 'h107b4, 'h107c4, 'h10a65, 'h107d4, 'h107e4, 'h10a66, 'h107f4, 'h10804, 'h10a67, 'h10814, 'h10824, 'h10a68, 'h103bc, 'h10834, 'h10844, 'h10a69, 'h10c64, 'h21f8e, 'h21f8f, 'h21f8d, 'h10854, 'h10864, 'h10a6a, 'h10874, 'h10884, 'h10a6b, 'h10894, 'h108a4, 'h10a6c, 'h108b4, 'h108c4, 'h10a6d, 'h108d4, 'h103bc, 'h106e4, 'h10a6e, 'h10c74, 'h106f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10704, 'h10a6f, 'h10714, 'h10724, 'h10a70, 'h10734, 'h10744, 'h10a71, 'h10754, 'h10764, 'h10a72, 'h10774, 'h10784, 'h10a73, 'h103bc, 'h10794, 'h10c74, 'h107a4, 'h10a74, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b4, 'h107c4, 'h10a75, 'h107d4, 'h107e4, 'h10a76, 'h107f4, 'h10804, 'h10a77, 'h10814, 'h10824, 'h10a78, 'h10834, 'h103bc, 'h10844, 'h10a79, 'h10c74, 'h10854, 'h21f8e, 'h21f8f, 'h21f8d, 'h10864, 'h10a7a, 'h10874, 'h10884, 'h10a7b, 'h10894, 'h108a4, 'h10a7c, 'h108b4, 'h108c4, 'h10a7d, 'h108d4, 'h106e4, 'h10a7e, 'h10c84, 'h103bc, 'h106f4, 'h10704, 'h10a7f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10714, 'h10724, 'h10a80, 'h10734, 'h10744, 'h10a81, 'h10754, 'h10764, 'h10a82, 'h10774, 'h10784, 'h10a83, 'h10794, 'h10c84, 'h103bc, 'h107a4, 'h10a84, 'h107b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c4, 'h10a85, 'h107d4, 'h107e4, 'h10a86, 'h107f4, 'h10804, 'h10a87, 'h10814, 'h10824, 'h10a88, 'h10834, 'h10844, 'h10a89, 'h10c84, 'h103bc, 'h10854, 'h10864, 'h10a8a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10874, 'h10884, 'h10a8b, 'h10894, 'h108a4, 'h10a8c, 'h108b4, 'h108c4, 'h10a8d, 'h108d4, 'h106e4, 'h10a8e, 'h10c94, 'h106f4, 'h103bc, 'h10704, 'h10a8f, 'h10714, 'h21f8e, 'h21f8f, 'h21f8d, 'h10724, 'h10a90, 'h10734, 'h10744, 'h10a91, 'h10754, 'h10764, 'h10a92, 'h10774, 'h10784, 'h10a93, 'h10794, 'h10c94, 'h107a4, 'h10a94, 'h103bc, 'h107b4, 'h107c4, 'h10a95, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d4, 'h107e4, 'h10a96, 'h107f4, 'h10804, 'h10a97, 'h10814, 'h10824, 'h10a98, 'h10834, 'h10844, 'h10a99, 'h10c94, 'h10854, 'h103bc, 'h10864, 'h10a9a, 'h10874, 'h21f8e, 'h21f8f, 'h21f8d, 'h10884, 'h10a9b, 'h10894, 'h108a4, 'h10a9c, 'h108b4, 'h108c4, 'h10a9d, 'h108d4, 'h106e4, 'h10a9e, 'h10ca4, 'h106f4, 'h10704, 'h10a9f, 'h103bc, 'h10714, 'h10724, 'h10aa0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10734, 'h10744, 'h10aa1, 'h10754, 'h10764, 'h10aa2, 'h10774, 'h10784, 'h10aa3, 'h10794, 'h10ca4, 'h107a4, 'h10aa4, 'h107b4, 'h103bc, 'h107c4, 'h10aa5, 'h107d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e4, 'h10aa6, 'h107f4, 'h10804, 'h10aa7, 'h10814, 'h10824, 'h10aa8, 'h10834, 'h10844, 'h10aa9, 'h10ca4, 'h10854, 'h10864, 'h10aaa, 'h103bc, 'h10874, 'h10884, 'h10aab, 'h21f8e, 'h21f8f, 'h21f8d, 'h10894, 'h108a4, 'h10aac, 'h108b4, 'h108c4, 'h10aad, 'h108d4, 'h106e4, 'h10aae, 'h10cb4, 'h106f4, 'h10704, 'h10aaf, 'h10714, 'h103bc, 'h10724, 'h10ab0, 'h10734, 'h21f8e, 'h21f8f, 'h21f8d, 'h10744, 'h10ab1, 'h10754, 'h10764, 'h10ab2, 'h10774, 'h10784, 'h10ab3, 'h10794, 'h10cb4, 'h107a4, 'h10ab4, 'h107b4, 'h107c4, 'h10ab5, 'h103bc, 'h107d4, 'h107e4, 'h10ab6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f4, 'h10804, 'h10ab7, 'h10814, 'h10824, 'h10ab8, 'h10834, 'h10844, 'h10ab9, 'h10cb4, 'h10854, 'h10864, 'h10aba, 'h10874, 'h103bc, 'h10884, 'h10abb, 'h10894, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a4, 'h10abc, 'h108b4, 'h108c4, 'h10abd, 'h108d4, 'h106e4, 'h10abe, 'h10cc4, 'h106f4, 'h10704, 'h10abf, 'h10714, 'h10724, 'h10ac0, 'h103bc, 'h10734, 'h10744, 'h10ac1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10754, 'h10764, 'h10ac2, 'h10774, 'h10784, 'h10ac3, 'h10794, 'h10cc4, 'h107a4, 'h10ac4, 'h107b4, 'h107c4, 'h10ac5, 'h107d4, 'h103bc, 'h107e4, 'h10ac6, 'h107f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10804, 'h10ac7, 'h10814, 'h10824, 'h10ac8, 'h10834, 'h10844, 'h10ac9, 'h10cc4, 'h10854, 'h10864, 'h10aca, 'h10874, 'h10884, 'h10acb, 'h103bc, 'h10894, 'h108a4, 'h10acc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b4, 'h108c4, 'h10acd, 'h108d4, 'h106e4, 'h10ace, 'h10cd4, 'h106f4, 'h10704, 'h10acf, 'h10714, 'h10724, 'h10ad0, 'h10734, 'h103bc, 'h10744, 'h10ad1, 'h10754, 'h21f8e, 'h21f8f, 'h21f8d, 'h10764, 'h10ad2, 'h10774, 'h10784, 'h10ad3, 'h10794, 'h10cd4, 'h107a4, 'h10ad4, 'h107b4, 'h107c4, 'h10ad5, 'h107d4, 'h107e4, 'h10ad6, 'h103bc, 'h107f4, 'h10804, 'h10ad7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10814, 'h10824, 'h10ad8, 'h10834, 'h10844, 'h10ad9, 'h10cd4, 'h10854, 'h10864, 'h10ada, 'h10874, 'h10884, 'h10adb, 'h10894, 'h103bc, 'h108a4, 'h10adc, 'h108b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c4, 'h10add, 'h108d4, 'h106e4, 'h108de, 'h10ae4, 'h106f4, 'h10704, 'h108df, 'h10714, 'h10724, 'h108e0, 'h10734, 'h10744, 'h108e1, 'h103bc, 'h10754, 'h10764, 'h108e2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10774, 'h10784, 'h108e3, 'h10794, 'h10ae4, 'h107a4, 'h108e4, 'h107b4, 'h107c4, 'h108e5, 'h107d4, 'h107e4, 'h108e6, 'h107f4, 'h103bc, 'h10804, 'h108e7, 'h10814, 'h21f8e, 'h21f8f, 'h21f8d, 'h10824, 'h108e8, 'h10834, 'h10844, 'h108e9, 'h10ae4, 'h10854, 'h10864, 'h108ea, 'h10874, 'h10884, 'h108eb, 'h10894, 'h108a4, 'h108ec, 'h103bc, 'h108b4, 'h108c4, 'h108ed, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d4, 'h106e4, 'h108ee, 'h10af4, 'h106f4, 'h10704, 'h108ef, 'h10714, 'h10724, 'h108f0, 'h10734, 'h10744, 'h108f1, 'h10754, 'h103bc, 'h10764, 'h108f2, 'h10774, 'h21f8e, 'h21f8f, 'h21f8d, 'h10784, 'h108f3, 'h10794, 'h10af4, 'h107a4, 'h108f4, 'h107b4, 'h107c4, 'h108f5, 'h107d4, 'h107e4, 'h108f6, 'h107f4, 'h10804, 'h108f7, 'h103bc, 'h10814, 'h10824, 'h108f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10834, 'h10844, 'h108f9, 'h10af4, 'h10854, 'h10864, 'h108fa, 'h10874, 'h10884, 'h108fb, 'h10894, 'h108a4, 'h108fc, 'h108b4, 'h103bc, 'h108c4, 'h108fd, 'h108d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h108fe, 'h10b04, 'h106f4, 'h10704, 'h108ff, 'h10714, 'h10724, 'h10900, 'h10734, 'h10744, 'h10901, 'h10754, 'h10764, 'h10902, 'h103bc, 'h10774, 'h10784, 'h10903, 'h21f8e, 'h21f8f, 'h21f8d, 'h10794, 'h10b04, 'h107a4, 'h10904, 'h107b4, 'h107c4, 'h10905, 'h107d4, 'h107e4, 'h10906, 'h107f4, 'h10804, 'h10907, 'h10814, 'h103bc, 'h10824, 'h10908, 'h10834, 'h21f8e, 'h21f8f, 'h21f8d, 'h10844, 'h10909, 'h10b04, 'h10854, 'h10864, 'h1090a, 'h10874, 'h10884, 'h1090b, 'h10894, 'h108a4, 'h1090c, 'h108b4, 'h108c4, 'h1090d, 'h103bc, 'h108d4, 'h106e4, 'h1090e, 'h10b14, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f4, 'h10704, 'h1090f, 'h10714, 'h10724, 'h10910, 'h10734, 'h10744, 'h10911, 'h10754, 'h10764, 'h10912, 'h10774, 'h103bc, 'h10784, 'h10913, 'h10794, 'h10b14, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a4, 'h10914, 'h107b4, 'h107c4, 'h10915, 'h107d4, 'h107e4, 'h10916, 'h107f4, 'h10804, 'h10917, 'h10814, 'h10824, 'h10918, 'h103bc, 'h10834, 'h10844, 'h10919, 'h10b14, 'h21f8e, 'h21f8f, 'h21f8d, 'h10854, 'h10864, 'h1091a, 'h10874, 'h10884, 'h1091b, 'h10894, 'h108a4, 'h1091c, 'h108b4, 'h108c4, 'h1091d, 'h108d4, 'h103bc, 'h106e4, 'h1091e, 'h10b24, 'h106f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10704, 'h1091f, 'h10714, 'h10724, 'h10920, 'h10734, 'h10744, 'h10921, 'h10754, 'h10764, 'h10922, 'h10774, 'h10784, 'h10923, 'h103bc, 'h10794, 'h10b24, 'h107a4, 'h10924, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b4, 'h107c4, 'h10925, 'h107d4, 'h107e4, 'h10926, 'h107f4, 'h10804, 'h10927, 'h10814, 'h10824, 'h10928, 'h10834, 'h103bc, 'h10844, 'h10929, 'h10b24, 'h10854, 'h21f8e, 'h21f8f, 'h21f8d, 'h10864, 'h1092a, 'h10874, 'h10884, 'h1092b, 'h10894, 'h108a4, 'h1092c, 'h108b4, 'h108c4, 'h1092d, 'h108d4, 'h106e4, 'h1092e, 'h10b34, 'h103bc, 'h106f4, 'h10704, 'h1092f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10714, 'h10724, 'h10930, 'h10734, 'h10744, 'h10931, 'h10754, 'h10764, 'h10932, 'h10774, 'h10784, 'h10933, 'h10794, 'h10b34, 'h103bc, 'h107a4, 'h10934, 'h107b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c4, 'h10935, 'h107d4, 'h107e4, 'h10936, 'h107f4, 'h10804, 'h10937, 'h10814, 'h10824, 'h10938, 'h10834, 'h10844, 'h10939, 'h10b34, 'h103bc, 'h10854, 'h10864, 'h1093a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10874, 'h10884, 'h1093b, 'h10894, 'h108a4, 'h1093c, 'h108b4, 'h108c4, 'h1093d, 'h108d4, 'h106e4, 'h1093e, 'h10b44, 'h106f4, 'h103bc, 'h10704, 'h1093f, 'h10714, 'h21f8e, 'h21f8f, 'h21f8d, 'h10724, 'h10940, 'h10734, 'h10744, 'h10941, 'h10754, 'h10764, 'h10942, 'h10774, 'h10784, 'h10943, 'h10794, 'h10b44, 'h107a4, 'h10944, 'h103bc, 'h107b4, 'h107c4, 'h10945, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d4, 'h107e4, 'h10946, 'h107f4, 'h10804, 'h10947, 'h10814, 'h10824, 'h10948, 'h10834, 'h10844, 'h10949, 'h10b44, 'h10854, 'h103bc, 'h10864, 'h1094a, 'h10874, 'h21f8e, 'h21f8f, 'h21f8d, 'h10884, 'h1094b, 'h10894, 'h108a4, 'h1094c, 'h108b4, 'h108c4, 'h1094d, 'h108d4, 'h106e4, 'h1094e, 'h10b54, 'h106f4, 'h10704, 'h1094f, 'h103bc, 'h10714, 'h10724, 'h10950, 'h21f8e, 'h21f8f, 'h21f8d, 'h10734, 'h10744, 'h10951, 'h10754, 'h10764, 'h10952, 'h10774, 'h10784, 'h10953, 'h10794, 'h10b54, 'h107a4, 'h10954, 'h107b4, 'h103bc, 'h107c4, 'h10955, 'h107d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e4, 'h10956, 'h107f4, 'h10804, 'h10957, 'h10814, 'h10824, 'h10958, 'h10834, 'h10844, 'h10959, 'h10b54, 'h10854, 'h10864, 'h1095a, 'h103bc, 'h10874, 'h10884, 'h1095b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10894, 'h108a4, 'h1095c, 'h108b4, 'h108c4, 'h1095d, 'h108d4, 'h106e4, 'h1095e, 'h10b64, 'h106f4, 'h10704, 'h1095f, 'h10714, 'h103bc, 'h10724, 'h10960, 'h10734, 'h21f8e, 'h21f8f, 'h21f8d, 'h10744, 'h10961, 'h10754, 'h10764, 'h10962, 'h10774, 'h10784, 'h10963, 'h10794, 'h10b64, 'h107a4, 'h10964, 'h107b4, 'h107c4, 'h10965, 'h103bc, 'h107d4, 'h107e4, 'h10966, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f4, 'h10804, 'h10967, 'h10814, 'h10824, 'h10968, 'h10834, 'h10844, 'h10969, 'h10b64, 'h10854, 'h10864, 'h1096a, 'h10874, 'h103bc, 'h10884, 'h1096b, 'h10894, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a4, 'h1096c, 'h108b4, 'h108c4, 'h1096d, 'h108d4, 'h106e4, 'h1096e, 'h10b74, 'h106f4, 'h10704, 'h1096f, 'h10714, 'h10724, 'h10970, 'h103bc, 'h10734, 'h10744, 'h10971, 'h21f8e, 'h21f8f, 'h21f8d, 'h10754, 'h10764, 'h10972, 'h10774, 'h10784, 'h10973, 'h10794, 'h10b74, 'h107a4, 'h10974, 'h107b4, 'h107c4, 'h10975, 'h107d4, 'h103bc, 'h107e4, 'h10976, 'h107f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10804, 'h10977, 'h10814, 'h10824, 'h10978, 'h10834, 'h10844, 'h10979, 'h10b74, 'h10854, 'h10864, 'h1097a, 'h10874, 'h10884, 'h1097b, 'h103bc, 'h10894, 'h108a4, 'h1097c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b4, 'h108c4, 'h1097d, 'h108d4, 'h106e4, 'h1097e, 'h10b84, 'h106f4, 'h10704, 'h1097f, 'h10714, 'h10724, 'h10980, 'h10734, 'h103bc, 'h10744, 'h10981, 'h10754, 'h21f8e, 'h21f8f, 'h21f8d, 'h10764, 'h10982, 'h10774, 'h10784, 'h10983, 'h10794, 'h10b84, 'h107a4, 'h10984, 'h107b4, 'h107c4, 'h10985, 'h107d4, 'h107e4, 'h10986, 'h103bc, 'h107f4, 'h10804, 'h10987, 'h21f8e, 'h21f8f, 'h21f8d, 'h10814, 'h10824, 'h10988, 'h10834, 'h10844, 'h10989, 'h10b84, 'h10854, 'h10864, 'h1098a, 'h10874, 'h10884, 'h1098b, 'h10894, 'h103bc, 'h108a4, 'h1098c, 'h108b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c4, 'h1098d, 'h108d4, 'h106e4, 'h1098e, 'h10b94, 'h106f4, 'h10704, 'h1098f, 'h10714, 'h10724, 'h10990, 'h10734, 'h10744, 'h10991, 'h103bc, 'h10754, 'h10764, 'h10992, 'h21f8e, 'h21f8f, 'h21f8d, 'h10774, 'h10784, 'h10993, 'h10794, 'h10b94, 'h107a4, 'h10994, 'h107b4, 'h107c4, 'h10995, 'h107d4, 'h107e4, 'h10996, 'h107f4, 'h103bc, 'h10804, 'h10997, 'h10814, 'h21f8e, 'h21f8f, 'h21f8d, 'h10824, 'h10998, 'h10834, 'h10844, 'h10999, 'h10b94, 'h10854, 'h10864, 'h1099a, 'h10874, 'h10884, 'h1099b, 'h10894, 'h108a4, 'h1099c, 'h103bc, 'h108b4, 'h108c4, 'h1099d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d4, 'h106e4, 'h1099e, 'h10ba4, 'h106f4, 'h10704, 'h1099f, 'h10714, 'h10724, 'h109a0, 'h10734, 'h10744, 'h109a1, 'h10754, 'h103bc, 'h10764, 'h109a2, 'h10774, 'h21f8e, 'h21f8f, 'h21f8d, 'h10784, 'h109a3, 'h10794, 'h10ba4, 'h107a4, 'h109a4, 'h107b4, 'h107c4, 'h109a5, 'h107d4, 'h107e4, 'h109a6, 'h107f4, 'h10804, 'h109a7, 'h103bc, 'h10814, 'h10824, 'h109a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10834, 'h10844, 'h109a9, 'h10ba4, 'h10854, 'h10864, 'h109aa, 'h10874, 'h10884, 'h109ab, 'h10894, 'h108a4, 'h109ac, 'h108b4, 'h103bc, 'h108c4, 'h109ad, 'h108d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h109ae, 'h10bb4, 'h106f4, 'h10704, 'h109af, 'h10714, 'h10724, 'h109b0, 'h10734, 'h10744, 'h109b1, 'h10754, 'h10764, 'h109b2, 'h103bc, 'h10774, 'h10784, 'h109b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10794, 'h10bb4, 'h107a4, 'h109b4, 'h107b4, 'h107c4, 'h109b5, 'h107d4, 'h107e4, 'h109b6, 'h107f4, 'h10804, 'h109b7, 'h10814, 'h103bc, 'h10824, 'h109b8, 'h10834, 'h21f8e, 'h21f8f, 'h21f8d, 'h10844, 'h109b9, 'h10bb4, 'h10854, 'h10864, 'h109ba, 'h10874, 'h10884, 'h109bb, 'h10894, 'h108a4, 'h109bc, 'h108b4, 'h108c4, 'h109bd, 'h103bc, 'h108d4, 'h106e4, 'h109be, 'h10bc4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f4, 'h10704, 'h109bf, 'h10714, 'h10724, 'h109c0, 'h10734, 'h10744, 'h109c1, 'h10754, 'h10764, 'h109c2, 'h10774, 'h103bc, 'h10784, 'h109c3, 'h10794, 'h10bc4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a4, 'h109c4, 'h107b4, 'h107c4, 'h109c5, 'h107d4, 'h107e4, 'h109c6, 'h107f4, 'h10804, 'h109c7, 'h10814, 'h10824, 'h109c8, 'h103bc, 'h10834, 'h10844, 'h109c9, 'h10bc4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10854, 'h10864, 'h109ca, 'h10874, 'h10884, 'h109cb, 'h10894, 'h108a4, 'h109cc, 'h108b4, 'h108c4, 'h109cd, 'h108d4, 'h103bc, 'h106e4, 'h109ce, 'h10bd4, 'h106f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10704, 'h109cf, 'h10714, 'h10724, 'h109d0, 'h10734, 'h10744, 'h109d1, 'h10754, 'h10764, 'h109d2, 'h10774, 'h10784, 'h109d3, 'h103bc, 'h10794, 'h10bd4, 'h107a4, 'h109d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b4, 'h107c4, 'h109d5, 'h107d4, 'h107e4, 'h109d6, 'h107f4, 'h10804, 'h109d7, 'h10814, 'h10824, 'h109d8, 'h10834, 'h103bc, 'h10844, 'h109d9, 'h10bd4, 'h10854, 'h21f8e, 'h21f8f, 'h21f8d, 'h10864, 'h109da, 'h10874, 'h10884, 'h109db, 'h10894, 'h108a4, 'h109dc, 'h108b4, 'h108c4, 'h109dd, 'h108d4, 'h106e4, 'h109de, 'h10be4, 'h103bc, 'h106f4, 'h10704, 'h109df, 'h21f8e, 'h21f8f, 'h21f8d, 'h10714, 'h10724, 'h109e0, 'h10734, 'h10744, 'h109e1, 'h10754, 'h10764, 'h109e2, 'h10774, 'h10784, 'h109e3, 'h10794, 'h10be4, 'h103bc, 'h107a4, 'h109e4, 'h107b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c4, 'h109e5, 'h107d4, 'h107e4, 'h109e6, 'h107f4, 'h10804, 'h109e7, 'h10814, 'h10824, 'h109e8, 'h10834, 'h10844, 'h109e9, 'h10be4, 'h103bc, 'h10854, 'h10864, 'h109ea, 'h21f8e, 'h21f8f, 'h21f8d, 'h10874, 'h10884, 'h109eb, 'h10894, 'h108a4, 'h109ec, 'h108b4, 'h108c4, 'h109ed, 'h108d4, 'h106e4, 'h109ee, 'h10bf4, 'h106f4, 'h103bc, 'h10704, 'h109ef, 'h10714, 'h21f8e, 'h21f8f, 'h21f8d, 'h10724, 'h109f0, 'h10734, 'h10744, 'h109f1, 'h10754, 'h10764, 'h109f2, 'h10774, 'h10784, 'h109f3, 'h10794, 'h10bf4, 'h107a4, 'h109f4, 'h103bc, 'h107b4, 'h107c4, 'h109f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d4, 'h107e4, 'h109f6, 'h107f4, 'h10804, 'h109f7, 'h10814, 'h10824, 'h109f8, 'h10834, 'h10844, 'h109f9, 'h10bf4, 'h10854, 'h103bc, 'h10864, 'h109fa, 'h10874, 'h21f8e, 'h21f8f, 'h21f8d, 'h10884, 'h109fb, 'h10894, 'h108a4, 'h109fc, 'h108b4, 'h108c4, 'h109fd, 'h108d4, 'h106e4, 'h109fe, 'h10c04, 'h106f4, 'h10704, 'h109ff, 'h103bc, 'h10714, 'h10724, 'h10a00, 'h21f8e, 'h21f8f, 'h21f8d, 'h10734, 'h10744, 'h10a01, 'h10754, 'h10764, 'h10a02, 'h10774, 'h10784, 'h10a03, 'h10794, 'h10c04, 'h107a4, 'h10a04, 'h107b4, 'h103bc, 'h107c4, 'h10a05, 'h107d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e4, 'h10a06, 'h107f4, 'h10804, 'h10a07, 'h10814, 'h10824, 'h10a08, 'h10834, 'h10844, 'h10a09, 'h10c04, 'h10854, 'h10864, 'h10a0a, 'h103bc, 'h10874, 'h10884, 'h10a0b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10894, 'h108a4, 'h10a0c, 'h108b4, 'h108c4, 'h10a0d, 'h108d4, 'h106e4, 'h10a0e, 'h10c14, 'h106f4, 'h10704, 'h10a0f, 'h10714, 'h103bc, 'h10724, 'h10a10, 'h10734, 'h21f8e, 'h21f8f, 'h21f8d, 'h10744, 'h10a11, 'h10754, 'h10764, 'h10a12, 'h10774, 'h10784, 'h10a13, 'h10794, 'h10c14, 'h107a4, 'h10a14, 'h107b4, 'h107c4, 'h10a15, 'h103bc, 'h107d4, 'h107e4, 'h10a16, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f4, 'h10804, 'h10a17, 'h10814, 'h10824, 'h10a18, 'h10834, 'h10844, 'h10a19, 'h10c14, 'h10854, 'h10864, 'h10a1a, 'h10874, 'h103bc, 'h10884, 'h10a1b, 'h10894, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a4, 'h10a1c, 'h108b4, 'h108c4, 'h10a1d, 'h108d4, 'h106e4, 'h10a1e, 'h10c24, 'h106f4, 'h10704, 'h10a1f, 'h10714, 'h10724, 'h10a20, 'h103bc, 'h10734, 'h10744, 'h10a21, 'h21f8e, 'h21f8f, 'h21f8d, 'h10754, 'h10764, 'h10a22, 'h10774, 'h10784, 'h10a23, 'h10794, 'h10c24, 'h107a4, 'h10a24, 'h107b4, 'h107c4, 'h10a25, 'h107d4, 'h103bc, 'h107e4, 'h10a26, 'h107f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10804, 'h10a27, 'h10814, 'h10824, 'h10a28, 'h10834, 'h10844, 'h10a29, 'h10c24, 'h10854, 'h10864, 'h10a2a, 'h10874, 'h10884, 'h10a2b, 'h103bc, 'h10894, 'h108a4, 'h10a2c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b4, 'h108c4, 'h10a2d, 'h108d4, 'h106e4, 'h10a2e, 'h10c34, 'h106f4, 'h10704, 'h10a2f, 'h10714, 'h10724, 'h10a30, 'h10734, 'h103bc, 'h10744, 'h10a31, 'h10754, 'h21f8e, 'h21f8f, 'h21f8d, 'h10764, 'h10a32, 'h10774, 'h10784, 'h10a33, 'h10794, 'h10c34, 'h107a4, 'h10a34, 'h107b4, 'h107c4, 'h10a35, 'h107d4, 'h107e4, 'h10a36, 'h103bc, 'h107f4, 'h10804, 'h10a37, 'h21f8e, 'h21f8f, 'h21f8d, 'h10814, 'h10824, 'h10a38, 'h10834, 'h10844, 'h10a39, 'h10c34, 'h10854, 'h10864, 'h10a3a, 'h10874, 'h10884, 'h10a3b, 'h10894, 'h103bc, 'h108a4, 'h10a3c, 'h108b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c4, 'h10a3d, 'h108d4, 'h106e4, 'h10a3e, 'h10c44, 'h106f4, 'h10704, 'h10a3f, 'h10714, 'h10724, 'h10a40, 'h10734, 'h10744, 'h10a41, 'h103bc, 'h10754, 'h10764, 'h10a42, 'h21f8e, 'h21f8f, 'h21f8d, 'h10774, 'h10784, 'h10a43, 'h10794, 'h10c44, 'h107a4, 'h10a44, 'h107b4, 'h107c4, 'h10a45, 'h107d4, 'h107e4, 'h10a46, 'h107f4, 'h103bc, 'h10804, 'h10a47, 'h10814, 'h21f8e, 'h21f8f, 'h21f8d, 'h10824, 'h10a48, 'h10834, 'h10844, 'h10a49, 'h10c44, 'h10854, 'h10864, 'h10a4a, 'h10874, 'h10884, 'h10a4b, 'h10894, 'h108a4, 'h10a4c, 'h103bc, 'h108b4, 'h108c4, 'h10a4d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d4, 'h106e4, 'h10a4e, 'h10c54, 'h106f4, 'h10704, 'h10a4f, 'h10714, 'h10724, 'h10a50, 'h10734, 'h10744, 'h10a51, 'h10754, 'h103bc, 'h10764, 'h10a52, 'h10774, 'h21f8e, 'h21f8f, 'h21f8d, 'h10784, 'h10a53, 'h10794, 'h10c54, 'h107a4, 'h10a54, 'h107b4, 'h107c4, 'h10a55, 'h107d4, 'h107e4, 'h10a56, 'h107f4, 'h10804, 'h10a57, 'h103bc, 'h10814, 'h10824, 'h10a58, 'h21f8e, 'h21f8f, 'h21f8d, 'h10834, 'h10844, 'h10a59, 'h10c54, 'h10854, 'h10864, 'h10a5a, 'h10874, 'h10884, 'h10a5b, 'h10894, 'h108a4, 'h10a5c, 'h108b4, 'h103bc, 'h108c4, 'h10a5d, 'h108d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h10a5e, 'h10c64, 'h106f4, 'h10704, 'h10a5f, 'h10714, 'h10724, 'h10a60, 'h10734, 'h10744, 'h10a61, 'h10754, 'h10764, 'h10a62, 'h103bc, 'h10774, 'h10784, 'h10a63, 'h21f8e, 'h21f8f, 'h21f8d, 'h10794, 'h10c64, 'h107a4, 'h10a64, 'h107b4, 'h107c4, 'h10a65, 'h107d4, 'h107e4, 'h10a66, 'h107f4, 'h10804, 'h10a67, 'h10814, 'h103bc, 'h10824, 'h10a68, 'h10834, 'h21f8e, 'h21f8f, 'h21f8d, 'h10844, 'h10a69, 'h10c64, 'h10854, 'h10864, 'h10a6a, 'h10874, 'h10884, 'h10a6b, 'h10894, 'h108a4, 'h10a6c, 'h108b4, 'h108c4, 'h10a6d, 'h103bc, 'h108d4, 'h106e4, 'h10a6e, 'h10c74, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f4, 'h10704, 'h10a6f, 'h10714, 'h10724, 'h10a70, 'h10734, 'h10744, 'h10a71, 'h10754, 'h10764, 'h10a72, 'h10774, 'h103bc, 'h10784, 'h10a73, 'h10794, 'h10c74, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a4, 'h10a74, 'h107b4, 'h107c4, 'h10a75, 'h107d4, 'h107e4, 'h10a76, 'h107f4, 'h10804, 'h10a77, 'h10814, 'h10824, 'h10a78, 'h103bc, 'h10834, 'h10844, 'h10a79, 'h10c74, 'h21f8e, 'h21f8f, 'h21f8d, 'h10854, 'h10864, 'h10a7a, 'h10874, 'h10884, 'h10a7b, 'h10894, 'h108a4, 'h10a7c, 'h108b4, 'h108c4, 'h10a7d, 'h108d4, 'h103bc, 'h106e4, 'h10a7e, 'h10c84, 'h106f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10704, 'h10a7f, 'h10714, 'h10724, 'h10a80, 'h10734, 'h10744, 'h10a81, 'h10754, 'h10764, 'h10a82, 'h10774, 'h10784, 'h10a83, 'h103bc, 'h10794, 'h10c84, 'h107a4, 'h10a84, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b4, 'h107c4, 'h10a85, 'h107d4, 'h107e4, 'h10a86, 'h107f4, 'h10804, 'h10a87, 'h10814, 'h10824, 'h10a88, 'h10834, 'h103bc, 'h10844, 'h10a89, 'h10c84, 'h10854, 'h21f8e, 'h21f8f, 'h21f8d, 'h10864, 'h10a8a, 'h10874, 'h10884, 'h10a8b, 'h10894, 'h108a4, 'h10a8c, 'h108b4, 'h108c4, 'h10a8d, 'h108d4, 'h106e4, 'h10a8e, 'h10c94, 'h103bc, 'h106f4, 'h10704, 'h10a8f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10714, 'h10724, 'h10a90, 'h10734, 'h10744, 'h10a91, 'h10754, 'h10764, 'h10a92, 'h10774, 'h10784, 'h10a93, 'h10794, 'h10c94, 'h103bc, 'h107a4, 'h10a94, 'h107b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c4, 'h10a95, 'h107d4, 'h107e4, 'h10a96, 'h107f4, 'h10804, 'h10a97, 'h10814, 'h10824, 'h10a98, 'h10834, 'h10844, 'h10a99, 'h10c94, 'h103bc, 'h10854, 'h10864, 'h10a9a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10874, 'h10884, 'h10a9b, 'h10894, 'h108a4, 'h10a9c, 'h108b4, 'h108c4, 'h10a9d, 'h108d4, 'h106e4, 'h10a9e, 'h10ca4, 'h106f4, 'h103bc, 'h10704, 'h10a9f, 'h10714, 'h21f8e, 'h21f8f, 'h21f8d, 'h10724, 'h10aa0, 'h10734, 'h10744, 'h10aa1, 'h10754, 'h10764, 'h10aa2, 'h10774, 'h10784, 'h10aa3, 'h10794, 'h10ca4, 'h107a4, 'h10aa4, 'h103bc, 'h107b4, 'h107c4, 'h10aa5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d4, 'h107e4, 'h10aa6, 'h107f4, 'h10804, 'h10aa7, 'h10814, 'h10824, 'h10aa8, 'h10834, 'h10844, 'h10aa9, 'h10ca4, 'h10854, 'h103bc, 'h10864, 'h10aaa, 'h10874, 'h21f8e, 'h21f8f, 'h21f8d, 'h10884, 'h10aab, 'h10894, 'h108a4, 'h10aac, 'h108b4, 'h108c4, 'h10aad, 'h108d4, 'h106e4, 'h10aae, 'h10cb4, 'h106f4, 'h10704, 'h10aaf, 'h103bc, 'h10714, 'h10724, 'h10ab0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10734, 'h10744, 'h10ab1, 'h10754, 'h10764, 'h10ab2, 'h10774, 'h10784, 'h10ab3, 'h10794, 'h10cb4, 'h107a4, 'h10ab4, 'h107b4, 'h103bc, 'h107c4, 'h10ab5, 'h107d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e4, 'h10ab6, 'h107f4, 'h10804, 'h10ab7, 'h10814, 'h10824, 'h10ab8, 'h10834, 'h10844, 'h10ab9, 'h10cb4, 'h10854, 'h10864, 'h10aba, 'h103bc, 'h10874, 'h10884, 'h10abb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10894, 'h108a4, 'h10abc, 'h108b4, 'h108c4, 'h10abd, 'h108d4, 'h106e4, 'h10abe, 'h10cc4, 'h106f4, 'h10704, 'h10abf, 'h10714, 'h103bc, 'h10724, 'h10ac0, 'h10734, 'h21f8e, 'h21f8f, 'h21f8d, 'h10744, 'h10ac1, 'h10754, 'h10764, 'h10ac2, 'h10774, 'h10784, 'h10ac3, 'h10794, 'h10cc4, 'h107a4, 'h10ac4, 'h107b4, 'h107c4, 'h10ac5, 'h103bc, 'h107d4, 'h107e4, 'h10ac6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f4, 'h10804, 'h10ac7, 'h10814, 'h10824, 'h10ac8, 'h10834, 'h10844, 'h10ac9, 'h10cc4, 'h10854, 'h10864, 'h10aca, 'h10874, 'h103bc, 'h10884, 'h10acb, 'h10894, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a4, 'h10acc, 'h108b4, 'h108c4, 'h10acd, 'h108d4, 'h106e4, 'h10ace, 'h10cd4, 'h106f4, 'h10704, 'h10acf, 'h10714, 'h10724, 'h10ad0, 'h103bc, 'h10734, 'h10744, 'h10ad1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10754, 'h10764, 'h10ad2, 'h10774, 'h10784, 'h10ad3, 'h10794, 'h10cd4, 'h107a4, 'h10ad4, 'h107b4, 'h107c4, 'h10ad5, 'h107d4, 'h103bc, 'h107e4, 'h10ad6, 'h107f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h10804, 'h10ad7, 'h10814, 'h10824, 'h10ad8, 'h10834, 'h10844, 'h10ad9, 'h10cd4, 'h10854, 'h10864, 'h10ada, 'h10874, 'h10884, 'h10adb, 'h103bc, 'h10894, 'h108a4, 'h10adc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b4, 'h108c4, 'h10add, 'h108d4, 'h106e5, 'h108de, 'h10ae5, 'h106f5, 'h10705, 'h108df, 'h10715, 'h10725, 'h108e0, 'h10735, 'h103bc, 'h10745, 'h108e1, 'h10755, 'h21f8e, 'h21f8f, 'h21f8d, 'h10765, 'h108e2, 'h10775, 'h10785, 'h108e3, 'h10795, 'h10ae5, 'h107a5, 'h108e4, 'h107b5, 'h107c5, 'h108e5, 'h107d5, 'h107e5, 'h108e6, 'h103bc, 'h107f5, 'h10805, 'h108e7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10815, 'h10825, 'h108e8, 'h10835, 'h10845, 'h108e9, 'h10ae5, 'h10855, 'h10865, 'h108ea, 'h10875, 'h10885, 'h108eb, 'h10895, 'h103bc, 'h108a5, 'h108ec, 'h108b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c5, 'h108ed, 'h108d5, 'h106e5, 'h108ee, 'h10af5, 'h106f5, 'h10705, 'h108ef, 'h10715, 'h10725, 'h108f0, 'h10735, 'h10745, 'h108f1, 'h103bc, 'h10755, 'h10765, 'h108f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10775, 'h10785, 'h108f3, 'h10795, 'h10af5, 'h107a5, 'h108f4, 'h107b5, 'h107c5, 'h108f5, 'h107d5, 'h107e5, 'h108f6, 'h107f5, 'h103bc, 'h10805, 'h108f7, 'h10815, 'h21f8e, 'h21f8f, 'h21f8d, 'h10825, 'h108f8, 'h10835, 'h10845, 'h108f9, 'h10af5, 'h10855, 'h10865, 'h108fa, 'h10875, 'h10885, 'h108fb, 'h10895, 'h108a5, 'h108fc, 'h103bc, 'h108b5, 'h108c5, 'h108fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d5, 'h106e5, 'h108fe, 'h10b05, 'h106f5, 'h10705, 'h108ff, 'h10715, 'h10725, 'h10900, 'h10735, 'h10745, 'h10901, 'h10755, 'h103bc, 'h10765, 'h10902, 'h10775, 'h21f8e, 'h21f8f, 'h21f8d, 'h10785, 'h10903, 'h10795, 'h10b05, 'h107a5, 'h10904, 'h107b5, 'h107c5, 'h10905, 'h107d5, 'h107e5, 'h10906, 'h107f5, 'h10805, 'h10907, 'h103bc, 'h10815, 'h10825, 'h10908, 'h21f8e, 'h21f8f, 'h21f8d, 'h10835, 'h10845, 'h10909, 'h10b05, 'h10855, 'h10865, 'h1090a, 'h10875, 'h10885, 'h1090b, 'h10895, 'h108a5, 'h1090c, 'h108b5, 'h103bc, 'h108c5, 'h1090d, 'h108d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1090e, 'h10b15, 'h106f5, 'h10705, 'h1090f, 'h10715, 'h10725, 'h10910, 'h10735, 'h10745, 'h10911, 'h10755, 'h10765, 'h10912, 'h103bc, 'h10775, 'h10785, 'h10913, 'h21f8e, 'h21f8f, 'h21f8d, 'h10795, 'h10b15, 'h107a5, 'h10914, 'h107b5, 'h107c5, 'h10915, 'h107d5, 'h107e5, 'h10916, 'h107f5, 'h10805, 'h10917, 'h10815, 'h103bc, 'h10825, 'h10918, 'h10835, 'h21f8e, 'h21f8f, 'h21f8d, 'h10845, 'h10919, 'h10b15, 'h10855, 'h10865, 'h1091a, 'h10875, 'h10885, 'h1091b, 'h10895, 'h108a5, 'h1091c, 'h108b5, 'h108c5, 'h1091d, 'h103bc, 'h108d5, 'h106e5, 'h1091e, 'h10b25, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f5, 'h10705, 'h1091f, 'h10715, 'h10725, 'h10920, 'h10735, 'h10745, 'h10921, 'h10755, 'h10765, 'h10922, 'h10775, 'h103bc, 'h10785, 'h10923, 'h10795, 'h10b25, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a5, 'h10924, 'h107b5, 'h107c5, 'h10925, 'h107d5, 'h107e5, 'h10926, 'h107f5, 'h10805, 'h10927, 'h10815, 'h10825, 'h10928, 'h103bc, 'h10835, 'h10845, 'h10929, 'h10b25, 'h21f8e, 'h21f8f, 'h21f8d, 'h10855, 'h10865, 'h1092a, 'h10875, 'h10885, 'h1092b, 'h10895, 'h108a5, 'h1092c, 'h108b5, 'h108c5, 'h1092d, 'h108d5, 'h103bc, 'h106e5, 'h1092e, 'h10b35, 'h106f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10705, 'h1092f, 'h10715, 'h10725, 'h10930, 'h10735, 'h10745, 'h10931, 'h10755, 'h10765, 'h10932, 'h10775, 'h10785, 'h10933, 'h103bc, 'h10795, 'h10b35, 'h107a5, 'h10934, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b5, 'h107c5, 'h10935, 'h107d5, 'h107e5, 'h10936, 'h107f5, 'h10805, 'h10937, 'h10815, 'h10825, 'h10938, 'h10835, 'h103bc, 'h10845, 'h10939, 'h10b35, 'h10855, 'h21f8e, 'h21f8f, 'h21f8d, 'h10865, 'h1093a, 'h10875, 'h10885, 'h1093b, 'h10895, 'h108a5, 'h1093c, 'h108b5, 'h108c5, 'h1093d, 'h108d5, 'h106e5, 'h1093e, 'h10b45, 'h103bc, 'h106f5, 'h10705, 'h1093f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10715, 'h10725, 'h10940, 'h10735, 'h10745, 'h10941, 'h10755, 'h10765, 'h10942, 'h10775, 'h10785, 'h10943, 'h10795, 'h10b45, 'h103bc, 'h107a5, 'h10944, 'h107b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c5, 'h10945, 'h107d5, 'h107e5, 'h10946, 'h107f5, 'h10805, 'h10947, 'h10815, 'h10825, 'h10948, 'h10835, 'h10845, 'h10949, 'h10b45, 'h103bc, 'h10855, 'h10865, 'h1094a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10875, 'h10885, 'h1094b, 'h10895, 'h108a5, 'h1094c, 'h108b5, 'h108c5, 'h1094d, 'h108d5, 'h106e5, 'h1094e, 'h10b55, 'h106f5, 'h103bc, 'h10705, 'h1094f, 'h10715, 'h21f8e, 'h21f8f, 'h21f8d, 'h10725, 'h10950, 'h10735, 'h10745, 'h10951, 'h10755, 'h10765, 'h10952, 'h10775, 'h10785, 'h10953, 'h10795, 'h10b55, 'h107a5, 'h10954, 'h103bc, 'h107b5, 'h107c5, 'h10955, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d5, 'h107e5, 'h10956, 'h107f5, 'h10805, 'h10957, 'h10815, 'h10825, 'h10958, 'h10835, 'h10845, 'h10959, 'h10b55, 'h10855, 'h103bc, 'h10865, 'h1095a, 'h10875, 'h21f8e, 'h21f8f, 'h21f8d, 'h10885, 'h1095b, 'h10895, 'h108a5, 'h1095c, 'h108b5, 'h108c5, 'h1095d, 'h108d5, 'h106e5, 'h1095e, 'h10b65, 'h106f5, 'h10705, 'h1095f, 'h103bc, 'h10715, 'h10725, 'h10960, 'h21f8e, 'h21f8f, 'h21f8d, 'h10735, 'h10745, 'h10961, 'h10755, 'h10765, 'h10962, 'h10775, 'h10785, 'h10963, 'h10795, 'h10b65, 'h107a5, 'h10964, 'h107b5, 'h103bc, 'h107c5, 'h10965, 'h107d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e5, 'h10966, 'h107f5, 'h10805, 'h10967, 'h10815, 'h10825, 'h10968, 'h10835, 'h10845, 'h10969, 'h10b65, 'h10855, 'h10865, 'h1096a, 'h103bc, 'h10875, 'h10885, 'h1096b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10895, 'h108a5, 'h1096c, 'h108b5, 'h108c5, 'h1096d, 'h108d5, 'h106e5, 'h1096e, 'h10b75, 'h106f5, 'h10705, 'h1096f, 'h10715, 'h103bc, 'h10725, 'h10970, 'h10735, 'h21f8e, 'h21f8f, 'h21f8d, 'h10745, 'h10971, 'h10755, 'h10765, 'h10972, 'h10775, 'h10785, 'h10973, 'h10795, 'h10b75, 'h107a5, 'h10974, 'h107b5, 'h107c5, 'h10975, 'h103bc, 'h107d5, 'h107e5, 'h10976, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f5, 'h10805, 'h10977, 'h10815, 'h10825, 'h10978, 'h10835, 'h10845, 'h10979, 'h10b75, 'h10855, 'h10865, 'h1097a, 'h10875, 'h103bc, 'h10885, 'h1097b, 'h10895, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a5, 'h1097c, 'h108b5, 'h108c5, 'h1097d, 'h108d5, 'h106e5, 'h1097e, 'h10b85, 'h106f5, 'h10705, 'h1097f, 'h10715, 'h10725, 'h10980, 'h103bc, 'h10735, 'h10745, 'h10981, 'h21f8e, 'h21f8f, 'h21f8d, 'h10755, 'h10765, 'h10982, 'h10775, 'h10785, 'h10983, 'h10795, 'h10b85, 'h107a5, 'h10984, 'h107b5, 'h107c5, 'h10985, 'h107d5, 'h103bc, 'h107e5, 'h10986, 'h107f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10805, 'h10987, 'h10815, 'h10825, 'h10988, 'h10835, 'h10845, 'h10989, 'h10b85, 'h10855, 'h10865, 'h1098a, 'h10875, 'h10885, 'h1098b, 'h103bc, 'h10895, 'h108a5, 'h1098c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b5, 'h108c5, 'h1098d, 'h108d5, 'h106e5, 'h1098e, 'h10b95, 'h106f5, 'h10705, 'h1098f, 'h10715, 'h10725, 'h10990, 'h10735, 'h103bc, 'h10745, 'h10991, 'h10755, 'h21f8e, 'h21f8f, 'h21f8d, 'h10765, 'h10992, 'h10775, 'h10785, 'h10993, 'h10795, 'h10b95, 'h107a5, 'h10994, 'h107b5, 'h107c5, 'h10995, 'h107d5, 'h107e5, 'h10996, 'h103bc, 'h107f5, 'h10805, 'h10997, 'h21f8e, 'h21f8f, 'h21f8d, 'h10815, 'h10825, 'h10998, 'h10835, 'h10845, 'h10999, 'h10b95, 'h10855, 'h10865, 'h1099a, 'h10875, 'h10885, 'h1099b, 'h10895, 'h103bc, 'h108a5, 'h1099c, 'h108b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c5, 'h1099d, 'h108d5, 'h106e5, 'h1099e, 'h10ba5, 'h106f5, 'h10705, 'h1099f, 'h10715, 'h10725, 'h109a0, 'h10735, 'h10745, 'h109a1, 'h103bc, 'h10755, 'h10765, 'h109a2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10775, 'h10785, 'h109a3, 'h10795, 'h10ba5, 'h107a5, 'h109a4, 'h107b5, 'h107c5, 'h109a5, 'h107d5, 'h107e5, 'h109a6, 'h107f5, 'h103bc, 'h10805, 'h109a7, 'h10815, 'h21f8e, 'h21f8f, 'h21f8d, 'h10825, 'h109a8, 'h10835, 'h10845, 'h109a9, 'h10ba5, 'h10855, 'h10865, 'h109aa, 'h10875, 'h10885, 'h109ab, 'h10895, 'h108a5, 'h109ac, 'h103bc, 'h108b5, 'h108c5, 'h109ad, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d5, 'h106e5, 'h109ae, 'h10bb5, 'h106f5, 'h10705, 'h109af, 'h10715, 'h10725, 'h109b0, 'h10735, 'h10745, 'h109b1, 'h10755, 'h103bc, 'h10765, 'h109b2, 'h10775, 'h21f8e, 'h21f8f, 'h21f8d, 'h10785, 'h109b3, 'h10795, 'h10bb5, 'h107a5, 'h109b4, 'h107b5, 'h107c5, 'h109b5, 'h107d5, 'h107e5, 'h109b6, 'h107f5, 'h10805, 'h109b7, 'h103bc, 'h10815, 'h10825, 'h109b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10835, 'h10845, 'h109b9, 'h10bb5, 'h10855, 'h10865, 'h109ba, 'h10875, 'h10885, 'h109bb, 'h10895, 'h108a5, 'h109bc, 'h108b5, 'h103bc, 'h108c5, 'h109bd, 'h108d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h109be, 'h10bc5, 'h106f5, 'h10705, 'h109bf, 'h10715, 'h10725, 'h109c0, 'h10735, 'h10745, 'h109c1, 'h10755, 'h10765, 'h109c2, 'h103bc, 'h10775, 'h10785, 'h109c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10795, 'h10bc5, 'h107a5, 'h109c4, 'h107b5, 'h107c5, 'h109c5, 'h107d5, 'h107e5, 'h109c6, 'h107f5, 'h10805, 'h109c7, 'h10815, 'h103bc, 'h10825, 'h109c8, 'h10835, 'h21f8e, 'h21f8f, 'h21f8d, 'h10845, 'h109c9, 'h10bc5, 'h10855, 'h10865, 'h109ca, 'h10875, 'h10885, 'h109cb, 'h10895, 'h108a5, 'h109cc, 'h108b5, 'h108c5, 'h109cd, 'h103bc, 'h108d5, 'h106e5, 'h109ce, 'h10bd5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f5, 'h10705, 'h109cf, 'h10715, 'h10725, 'h109d0, 'h10735, 'h10745, 'h109d1, 'h10755, 'h10765, 'h109d2, 'h10775, 'h103bc, 'h10785, 'h109d3, 'h10795, 'h10bd5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a5, 'h109d4, 'h107b5, 'h107c5, 'h109d5, 'h107d5, 'h107e5, 'h109d6, 'h107f5, 'h10805, 'h109d7, 'h10815, 'h10825, 'h109d8, 'h103bc, 'h10835, 'h10845, 'h109d9, 'h10bd5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10855, 'h10865, 'h109da, 'h10875, 'h10885, 'h109db, 'h10895, 'h108a5, 'h109dc, 'h108b5, 'h108c5, 'h109dd, 'h108d5, 'h103bc, 'h106e5, 'h109de, 'h10be5, 'h106f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10705, 'h109df, 'h10715, 'h10725, 'h109e0, 'h10735, 'h10745, 'h109e1, 'h10755, 'h10765, 'h109e2, 'h10775, 'h10785, 'h109e3, 'h103bc, 'h10795, 'h10be5, 'h107a5, 'h109e4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b5, 'h107c5, 'h109e5, 'h107d5, 'h107e5, 'h109e6, 'h107f5, 'h10805, 'h109e7, 'h10815, 'h10825, 'h109e8, 'h10835, 'h103bc, 'h10845, 'h109e9, 'h10be5, 'h10855, 'h21f8e, 'h21f8f, 'h21f8d, 'h10865, 'h109ea, 'h10875, 'h10885, 'h109eb, 'h10895, 'h108a5, 'h109ec, 'h108b5, 'h108c5, 'h109ed, 'h108d5, 'h106e5, 'h109ee, 'h10bf5, 'h103bc, 'h106f5, 'h10705, 'h109ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h10715, 'h10725, 'h109f0, 'h10735, 'h10745, 'h109f1, 'h10755, 'h10765, 'h109f2, 'h10775, 'h10785, 'h109f3, 'h10795, 'h10bf5, 'h103bc, 'h107a5, 'h109f4, 'h107b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c5, 'h109f5, 'h107d5, 'h107e5, 'h109f6, 'h107f5, 'h10805, 'h109f7, 'h10815, 'h10825, 'h109f8, 'h10835, 'h10845, 'h109f9, 'h10bf5, 'h103bc, 'h10855, 'h10865, 'h109fa, 'h21f8e, 'h21f8f, 'h21f8d, 'h10875, 'h10885, 'h109fb, 'h10895, 'h108a5, 'h109fc, 'h108b5, 'h108c5, 'h109fd, 'h108d5, 'h106e5, 'h109fe, 'h10c05, 'h106f5, 'h103bc, 'h10705, 'h109ff, 'h10715, 'h21f8e, 'h21f8f, 'h21f8d, 'h10725, 'h10a00, 'h10735, 'h10745, 'h10a01, 'h10755, 'h10765, 'h10a02, 'h10775, 'h10785, 'h10a03, 'h10795, 'h10c05, 'h107a5, 'h10a04, 'h103bc, 'h107b5, 'h107c5, 'h10a05, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d5, 'h107e5, 'h10a06, 'h107f5, 'h10805, 'h10a07, 'h10815, 'h10825, 'h10a08, 'h10835, 'h10845, 'h10a09, 'h10c05, 'h10855, 'h103bc, 'h10865, 'h10a0a, 'h10875, 'h21f8e, 'h21f8f, 'h21f8d, 'h10885, 'h10a0b, 'h10895, 'h108a5, 'h10a0c, 'h108b5, 'h108c5, 'h10a0d, 'h108d5, 'h106e5, 'h10a0e, 'h10c15, 'h106f5, 'h10705, 'h10a0f, 'h103bc, 'h10715, 'h10725, 'h10a10, 'h21f8e, 'h21f8f, 'h21f8d, 'h10735, 'h10745, 'h10a11, 'h10755, 'h10765, 'h10a12, 'h10775, 'h10785, 'h10a13, 'h10795, 'h10c15, 'h107a5, 'h10a14, 'h107b5, 'h103bc, 'h107c5, 'h10a15, 'h107d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e5, 'h10a16, 'h107f5, 'h10805, 'h10a17, 'h10815, 'h10825, 'h10a18, 'h10835, 'h10845, 'h10a19, 'h10c15, 'h10855, 'h10865, 'h10a1a, 'h103bc, 'h10875, 'h10885, 'h10a1b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10895, 'h108a5, 'h10a1c, 'h108b5, 'h108c5, 'h10a1d, 'h108d5, 'h106e5, 'h10a1e, 'h10c25, 'h106f5, 'h10705, 'h10a1f, 'h10715, 'h103bc, 'h10725, 'h10a20, 'h10735, 'h21f8e, 'h21f8f, 'h21f8d, 'h10745, 'h10a21, 'h10755, 'h10765, 'h10a22, 'h10775, 'h10785, 'h10a23, 'h10795, 'h10c25, 'h107a5, 'h10a24, 'h107b5, 'h107c5, 'h10a25, 'h103bc, 'h107d5, 'h107e5, 'h10a26, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f5, 'h10805, 'h10a27, 'h10815, 'h10825, 'h10a28, 'h10835, 'h10845, 'h10a29, 'h10c25, 'h10855, 'h10865, 'h10a2a, 'h10875, 'h103bc, 'h10885, 'h10a2b, 'h10895, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a5, 'h10a2c, 'h108b5, 'h108c5, 'h10a2d, 'h108d5, 'h106e5, 'h10a2e, 'h10c35, 'h106f5, 'h10705, 'h10a2f, 'h10715, 'h10725, 'h10a30, 'h103bc, 'h10735, 'h10745, 'h10a31, 'h21f8e, 'h21f8f, 'h21f8d, 'h10755, 'h10765, 'h10a32, 'h10775, 'h10785, 'h10a33, 'h10795, 'h10c35, 'h107a5, 'h10a34, 'h107b5, 'h107c5, 'h10a35, 'h107d5, 'h103bc, 'h107e5, 'h10a36, 'h107f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10805, 'h10a37, 'h10815, 'h10825, 'h10a38, 'h10835, 'h10845, 'h10a39, 'h10c35, 'h10855, 'h10865, 'h10a3a, 'h10875, 'h10885, 'h10a3b, 'h103bc, 'h10895, 'h108a5, 'h10a3c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b5, 'h108c5, 'h10a3d, 'h108d5, 'h106e5, 'h10a3e, 'h10c45, 'h106f5, 'h10705, 'h10a3f, 'h10715, 'h10725, 'h10a40, 'h10735, 'h103bc, 'h10745, 'h10a41, 'h10755, 'h21f8e, 'h21f8f, 'h21f8d, 'h10765, 'h10a42, 'h10775, 'h10785, 'h10a43, 'h10795, 'h10c45, 'h107a5, 'h10a44, 'h107b5, 'h107c5, 'h10a45, 'h107d5, 'h107e5, 'h10a46, 'h103bc, 'h107f5, 'h10805, 'h10a47, 'h21f8e, 'h21f8f, 'h21f8d, 'h10815, 'h10825, 'h10a48, 'h10835, 'h10845, 'h10a49, 'h10c45, 'h10855, 'h10865, 'h10a4a, 'h10875, 'h10885, 'h10a4b, 'h10895, 'h103bc, 'h108a5, 'h10a4c, 'h108b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c5, 'h10a4d, 'h108d5, 'h106e5, 'h10a4e, 'h10c55, 'h106f5, 'h10705, 'h10a4f, 'h10715, 'h10725, 'h10a50, 'h10735, 'h10745, 'h10a51, 'h103bc, 'h10755, 'h10765, 'h10a52, 'h21f8e, 'h21f8f, 'h21f8d, 'h10775, 'h10785, 'h10a53, 'h10795, 'h10c55, 'h107a5, 'h10a54, 'h107b5, 'h107c5, 'h10a55, 'h107d5, 'h107e5, 'h10a56, 'h107f5, 'h103bc, 'h10805, 'h10a57, 'h10815, 'h21f8e, 'h21f8f, 'h21f8d, 'h10825, 'h10a58, 'h10835, 'h10845, 'h10a59, 'h10c55, 'h10855, 'h10865, 'h10a5a, 'h10875, 'h10885, 'h10a5b, 'h10895, 'h108a5, 'h10a5c, 'h103bc, 'h108b5, 'h108c5, 'h10a5d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d5, 'h106e5, 'h10a5e, 'h10c65, 'h106f5, 'h10705, 'h10a5f, 'h10715, 'h10725, 'h10a60, 'h10735, 'h10745, 'h10a61, 'h10755, 'h103bc, 'h10765, 'h10a62, 'h10775, 'h21f8e, 'h21f8f, 'h21f8d, 'h10785, 'h10a63, 'h10795, 'h10c65, 'h107a5, 'h10a64, 'h107b5, 'h107c5, 'h10a65, 'h107d5, 'h107e5, 'h10a66, 'h107f5, 'h10805, 'h10a67, 'h103bc, 'h10815, 'h10825, 'h10a68, 'h21f8e, 'h21f8f, 'h21f8d, 'h10835, 'h10845, 'h10a69, 'h10c65, 'h10855, 'h10865, 'h10a6a, 'h10875, 'h10885, 'h10a6b, 'h10895, 'h108a5, 'h10a6c, 'h108b5, 'h103bc, 'h108c5, 'h10a6d, 'h108d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h10a6e, 'h10c75, 'h106f5, 'h10705, 'h10a6f, 'h10715, 'h10725, 'h10a70, 'h10735, 'h10745, 'h10a71, 'h10755, 'h10765, 'h10a72, 'h103bc, 'h10775, 'h10785, 'h10a73, 'h21f8e, 'h21f8f, 'h21f8d, 'h10795, 'h10c75, 'h107a5, 'h10a74, 'h107b5, 'h107c5, 'h10a75, 'h107d5, 'h107e5, 'h10a76, 'h107f5, 'h10805, 'h10a77, 'h10815, 'h103bc, 'h10825, 'h10a78, 'h10835, 'h21f8e, 'h21f8f, 'h21f8d, 'h10845, 'h10a79, 'h10c75, 'h10855, 'h10865, 'h10a7a, 'h10875, 'h10885, 'h10a7b, 'h10895, 'h108a5, 'h10a7c, 'h108b5, 'h108c5, 'h10a7d, 'h103bc, 'h108d5, 'h106e5, 'h10a7e, 'h10c85, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f5, 'h10705, 'h10a7f, 'h10715, 'h10725, 'h10a80, 'h10735, 'h10745, 'h10a81, 'h10755, 'h10765, 'h10a82, 'h10775, 'h103bc, 'h10785, 'h10a83, 'h10795, 'h10c85, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a5, 'h10a84, 'h107b5, 'h107c5, 'h10a85, 'h107d5, 'h107e5, 'h10a86, 'h107f5, 'h10805, 'h10a87, 'h10815, 'h10825, 'h10a88, 'h103bc, 'h10835, 'h10845, 'h10a89, 'h10c85, 'h21f8e, 'h21f8f, 'h21f8d, 'h10855, 'h10865, 'h10a8a, 'h10875, 'h10885, 'h10a8b, 'h10895, 'h108a5, 'h10a8c, 'h108b5, 'h108c5, 'h10a8d, 'h108d5, 'h103bc, 'h106e5, 'h10a8e, 'h10c95, 'h106f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10705, 'h10a8f, 'h10715, 'h10725, 'h10a90, 'h10735, 'h10745, 'h10a91, 'h10755, 'h10765, 'h10a92, 'h10775, 'h10785, 'h10a93, 'h103bc, 'h10795, 'h10c95, 'h107a5, 'h10a94, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b5, 'h107c5, 'h10a95, 'h107d5, 'h107e5, 'h10a96, 'h107f5, 'h10805, 'h10a97, 'h10815, 'h10825, 'h10a98, 'h10835, 'h103bc, 'h10845, 'h10a99, 'h10c95, 'h10855, 'h21f8e, 'h21f8f, 'h21f8d, 'h10865, 'h10a9a, 'h10875, 'h10885, 'h10a9b, 'h10895, 'h108a5, 'h10a9c, 'h108b5, 'h108c5, 'h10a9d, 'h108d5, 'h106e5, 'h10a9e, 'h10ca5, 'h103bc, 'h106f5, 'h10705, 'h10a9f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10715, 'h10725, 'h10aa0, 'h10735, 'h10745, 'h10aa1, 'h10755, 'h10765, 'h10aa2, 'h10775, 'h10785, 'h10aa3, 'h10795, 'h10ca5, 'h103bc, 'h107a5, 'h10aa4, 'h107b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c5, 'h10aa5, 'h107d5, 'h107e5, 'h10aa6, 'h107f5, 'h10805, 'h10aa7, 'h10815, 'h10825, 'h10aa8, 'h10835, 'h10845, 'h10aa9, 'h10ca5, 'h103bc, 'h10855, 'h10865, 'h10aaa, 'h21f8e, 'h21f8f, 'h21f8d, 'h10875, 'h10885, 'h10aab, 'h10895, 'h108a5, 'h10aac, 'h108b5, 'h108c5, 'h10aad, 'h108d5, 'h106e5, 'h10aae, 'h10cb5, 'h106f5, 'h103bc, 'h10705, 'h10aaf, 'h10715, 'h21f8e, 'h21f8f, 'h21f8d, 'h10725, 'h10ab0, 'h10735, 'h10745, 'h10ab1, 'h10755, 'h10765, 'h10ab2, 'h10775, 'h10785, 'h10ab3, 'h10795, 'h10cb5, 'h107a5, 'h10ab4, 'h103bc, 'h107b5, 'h107c5, 'h10ab5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d5, 'h107e5, 'h10ab6, 'h107f5, 'h10805, 'h10ab7, 'h10815, 'h10825, 'h10ab8, 'h10835, 'h10845, 'h10ab9, 'h10cb5, 'h10855, 'h103bc, 'h10865, 'h10aba, 'h10875, 'h21f8e, 'h21f8f, 'h21f8d, 'h10885, 'h10abb, 'h10895, 'h108a5, 'h10abc, 'h108b5, 'h108c5, 'h10abd, 'h108d5, 'h106e5, 'h10abe, 'h10cc5, 'h106f5, 'h10705, 'h10abf, 'h103bc, 'h10715, 'h10725, 'h10ac0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10735, 'h10745, 'h10ac1, 'h10755, 'h10765, 'h10ac2, 'h10775, 'h10785, 'h10ac3, 'h10795, 'h10cc5, 'h107a5, 'h10ac4, 'h107b5, 'h103bc, 'h107c5, 'h10ac5, 'h107d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e5, 'h10ac6, 'h107f5, 'h10805, 'h10ac7, 'h10815, 'h10825, 'h10ac8, 'h10835, 'h10845, 'h10ac9, 'h10cc5, 'h10855, 'h10865, 'h10aca, 'h103bc, 'h10875, 'h10885, 'h10acb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10895, 'h108a5, 'h10acc, 'h108b5, 'h108c5, 'h10acd, 'h108d5, 'h106e5, 'h10ace, 'h10cd5, 'h106f5, 'h10705, 'h10acf, 'h10715, 'h103bc, 'h10725, 'h10ad0, 'h10735, 'h21f8e, 'h21f8f, 'h21f8d, 'h10745, 'h10ad1, 'h10755, 'h10765, 'h10ad2, 'h10775, 'h10785, 'h10ad3, 'h10795, 'h10cd5, 'h107a5, 'h10ad4, 'h107b5, 'h107c5, 'h10ad5, 'h103bc, 'h107d5, 'h107e5, 'h10ad6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f5, 'h10805, 'h10ad7, 'h10815, 'h10825, 'h10ad8, 'h10835, 'h10845, 'h10ad9, 'h10cd5, 'h10855, 'h10865, 'h10ada, 'h10875, 'h103bc, 'h10885, 'h10adb, 'h10895, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a5, 'h10adc, 'h108b5, 'h108c5, 'h10add, 'h108d5, 'h106e5, 'h108de, 'h10ae5, 'h106f5, 'h10705, 'h108df, 'h10715, 'h10725, 'h108e0, 'h103bc, 'h10735, 'h10745, 'h108e1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10755, 'h10765, 'h108e2, 'h10775, 'h10785, 'h108e3, 'h10795, 'h10ae5, 'h107a5, 'h108e4, 'h107b5, 'h107c5, 'h108e5, 'h107d5, 'h103bc, 'h107e5, 'h108e6, 'h107f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10805, 'h108e7, 'h10815, 'h10825, 'h108e8, 'h10835, 'h10845, 'h108e9, 'h10ae5, 'h10855, 'h10865, 'h108ea, 'h10875, 'h10885, 'h108eb, 'h103bc, 'h10895, 'h108a5, 'h108ec, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b5, 'h108c5, 'h108ed, 'h108d5, 'h106e5, 'h108ee, 'h10af5, 'h106f5, 'h10705, 'h108ef, 'h10715, 'h10725, 'h108f0, 'h10735, 'h103bc, 'h10745, 'h108f1, 'h10755, 'h21f8e, 'h21f8f, 'h21f8d, 'h10765, 'h108f2, 'h10775, 'h10785, 'h108f3, 'h10795, 'h10af5, 'h107a5, 'h108f4, 'h107b5, 'h107c5, 'h108f5, 'h107d5, 'h107e5, 'h108f6, 'h103bc, 'h107f5, 'h10805, 'h108f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10815, 'h10825, 'h108f8, 'h10835, 'h10845, 'h108f9, 'h10af5, 'h10855, 'h10865, 'h108fa, 'h10875, 'h10885, 'h108fb, 'h10895, 'h103bc, 'h108a5, 'h108fc, 'h108b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c5, 'h108fd, 'h108d5, 'h106e5, 'h108fe, 'h10b05, 'h106f5, 'h10705, 'h108ff, 'h10715, 'h10725, 'h10900, 'h10735, 'h10745, 'h10901, 'h103bc, 'h10755, 'h10765, 'h10902, 'h21f8e, 'h21f8f, 'h21f8d, 'h10775, 'h10785, 'h10903, 'h10795, 'h10b05, 'h107a5, 'h10904, 'h107b5, 'h107c5, 'h10905, 'h107d5, 'h107e5, 'h10906, 'h107f5, 'h103bc, 'h10805, 'h10907, 'h10815, 'h21f8e, 'h21f8f, 'h21f8d, 'h10825, 'h10908, 'h10835, 'h10845, 'h10909, 'h10b05, 'h10855, 'h10865, 'h1090a, 'h10875, 'h10885, 'h1090b, 'h10895, 'h108a5, 'h1090c, 'h103bc, 'h108b5, 'h108c5, 'h1090d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d5, 'h106e5, 'h1090e, 'h10b15, 'h106f5, 'h10705, 'h1090f, 'h10715, 'h10725, 'h10910, 'h10735, 'h10745, 'h10911, 'h10755, 'h103bc, 'h10765, 'h10912, 'h10775, 'h21f8e, 'h21f8f, 'h21f8d, 'h10785, 'h10913, 'h10795, 'h10b15, 'h107a5, 'h10914, 'h107b5, 'h107c5, 'h10915, 'h107d5, 'h107e5, 'h10916, 'h107f5, 'h10805, 'h10917, 'h103bc, 'h10815, 'h10825, 'h10918, 'h21f8e, 'h21f8f, 'h21f8d, 'h10835, 'h10845, 'h10919, 'h10b15, 'h10855, 'h10865, 'h1091a, 'h10875, 'h10885, 'h1091b, 'h10895, 'h108a5, 'h1091c, 'h108b5, 'h103bc, 'h108c5, 'h1091d, 'h108d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1091e, 'h10b25, 'h106f5, 'h10705, 'h1091f, 'h10715, 'h10725, 'h10920, 'h10735, 'h10745, 'h10921, 'h10755, 'h10765, 'h10922, 'h103bc, 'h10775, 'h10785, 'h10923, 'h21f8e, 'h21f8f, 'h21f8d, 'h10795, 'h10b25, 'h107a5, 'h10924, 'h107b5, 'h107c5, 'h10925, 'h107d5, 'h107e5, 'h10926, 'h107f5, 'h10805, 'h10927, 'h10815, 'h103bc, 'h10825, 'h10928, 'h10835, 'h21f8e, 'h21f8f, 'h21f8d, 'h10845, 'h10929, 'h10b25, 'h10855, 'h10865, 'h1092a, 'h10875, 'h10885, 'h1092b, 'h10895, 'h108a5, 'h1092c, 'h108b5, 'h108c5, 'h1092d, 'h103bc, 'h108d5, 'h106e5, 'h1092e, 'h10b35, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f5, 'h10705, 'h1092f, 'h10715, 'h10725, 'h10930, 'h10735, 'h10745, 'h10931, 'h10755, 'h10765, 'h10932, 'h10775, 'h103bc, 'h10785, 'h10933, 'h10795, 'h10b35, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a5, 'h10934, 'h107b5, 'h107c5, 'h10935, 'h107d5, 'h107e5, 'h10936, 'h107f5, 'h10805, 'h10937, 'h10815, 'h10825, 'h10938, 'h103bc, 'h10835, 'h10845, 'h10939, 'h10b35, 'h21f8e, 'h21f8f, 'h21f8d, 'h10855, 'h10865, 'h1093a, 'h10875, 'h10885, 'h1093b, 'h10895, 'h108a5, 'h1093c, 'h108b5, 'h108c5, 'h1093d, 'h108d5, 'h103bc, 'h106e5, 'h1093e, 'h10b45, 'h106f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10705, 'h1093f, 'h10715, 'h10725, 'h10940, 'h10735, 'h10745, 'h10941, 'h10755, 'h10765, 'h10942, 'h10775, 'h10785, 'h10943, 'h103bc, 'h10795, 'h10b45, 'h107a5, 'h10944, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b5, 'h107c5, 'h10945, 'h107d5, 'h107e5, 'h10946, 'h107f5, 'h10805, 'h10947, 'h10815, 'h10825, 'h10948, 'h10835, 'h103bc, 'h10845, 'h10949, 'h10b45, 'h10855, 'h21f8e, 'h21f8f, 'h21f8d, 'h10865, 'h1094a, 'h10875, 'h10885, 'h1094b, 'h10895, 'h108a5, 'h1094c, 'h108b5, 'h108c5, 'h1094d, 'h108d5, 'h106e5, 'h1094e, 'h10b55, 'h103bc, 'h106f5, 'h10705, 'h1094f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10715, 'h10725, 'h10950, 'h10735, 'h10745, 'h10951, 'h10755, 'h10765, 'h10952, 'h10775, 'h10785, 'h10953, 'h10795, 'h10b55, 'h103bc, 'h107a5, 'h10954, 'h107b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c5, 'h10955, 'h107d5, 'h107e5, 'h10956, 'h107f5, 'h10805, 'h10957, 'h10815, 'h10825, 'h10958, 'h10835, 'h10845, 'h10959, 'h10b55, 'h103bc, 'h10855, 'h10865, 'h1095a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10875, 'h10885, 'h1095b, 'h10895, 'h108a5, 'h1095c, 'h108b5, 'h108c5, 'h1095d, 'h108d5, 'h106e5, 'h1095e, 'h10b65, 'h106f5, 'h103bc, 'h10705, 'h1095f, 'h10715, 'h21f8e, 'h21f8f, 'h21f8d, 'h10725, 'h10960, 'h10735, 'h10745, 'h10961, 'h10755, 'h10765, 'h10962, 'h10775, 'h10785, 'h10963, 'h10795, 'h10b65, 'h107a5, 'h10964, 'h103bc, 'h107b5, 'h107c5, 'h10965, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d5, 'h107e5, 'h10966, 'h107f5, 'h10805, 'h10967, 'h10815, 'h10825, 'h10968, 'h10835, 'h10845, 'h10969, 'h10b65, 'h10855, 'h103bc, 'h10865, 'h1096a, 'h10875, 'h21f8e, 'h21f8f, 'h21f8d, 'h10885, 'h1096b, 'h10895, 'h108a5, 'h1096c, 'h108b5, 'h108c5, 'h1096d, 'h108d5, 'h106e5, 'h1096e, 'h10b75, 'h106f5, 'h10705, 'h1096f, 'h103bc, 'h10715, 'h10725, 'h10970, 'h21f8e, 'h21f8f, 'h21f8d, 'h10735, 'h10745, 'h10971, 'h10755, 'h10765, 'h10972, 'h10775, 'h10785, 'h10973, 'h10795, 'h10b75, 'h107a5, 'h10974, 'h107b5, 'h103bc, 'h107c5, 'h10975, 'h107d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e5, 'h10976, 'h107f5, 'h10805, 'h10977, 'h10815, 'h10825, 'h10978, 'h10835, 'h10845, 'h10979, 'h10b75, 'h10855, 'h10865, 'h1097a, 'h103bc, 'h10875, 'h10885, 'h1097b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10895, 'h108a5, 'h1097c, 'h108b5, 'h108c5, 'h1097d, 'h108d5, 'h106e5, 'h1097e, 'h10b85, 'h106f5, 'h10705, 'h1097f, 'h10715, 'h103bc, 'h10725, 'h10980, 'h10735, 'h21f8e, 'h21f8f, 'h21f8d, 'h10745, 'h10981, 'h10755, 'h10765, 'h10982, 'h10775, 'h10785, 'h10983, 'h10795, 'h10b85, 'h107a5, 'h10984, 'h107b5, 'h107c5, 'h10985, 'h103bc, 'h107d5, 'h107e5, 'h10986, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f5, 'h10805, 'h10987, 'h10815, 'h10825, 'h10988, 'h10835, 'h10845, 'h10989, 'h10b85, 'h10855, 'h10865, 'h1098a, 'h10875, 'h103bc, 'h10885, 'h1098b, 'h10895, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a5, 'h1098c, 'h108b5, 'h108c5, 'h1098d, 'h108d5, 'h106e5, 'h1098e, 'h10b95, 'h106f5, 'h10705, 'h1098f, 'h10715, 'h10725, 'h10990, 'h103bc, 'h10735, 'h10745, 'h10991, 'h21f8e, 'h21f8f, 'h21f8d, 'h10755, 'h10765, 'h10992, 'h10775, 'h10785, 'h10993, 'h10795, 'h10b95, 'h107a5, 'h10994, 'h107b5, 'h107c5, 'h10995, 'h107d5, 'h103bc, 'h107e5, 'h10996, 'h107f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10805, 'h10997, 'h10815, 'h10825, 'h10998, 'h10835, 'h10845, 'h10999, 'h10b95, 'h10855, 'h10865, 'h1099a, 'h10875, 'h10885, 'h1099b, 'h103bc, 'h10895, 'h108a5, 'h1099c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b5, 'h108c5, 'h1099d, 'h108d5, 'h106e5, 'h1099e, 'h10ba5, 'h106f5, 'h10705, 'h1099f, 'h10715, 'h10725, 'h109a0, 'h10735, 'h103bc, 'h10745, 'h109a1, 'h10755, 'h21f8e, 'h21f8f, 'h21f8d, 'h10765, 'h109a2, 'h10775, 'h10785, 'h109a3, 'h10795, 'h10ba5, 'h107a5, 'h109a4, 'h107b5, 'h107c5, 'h109a5, 'h107d5, 'h107e5, 'h109a6, 'h103bc, 'h107f5, 'h10805, 'h109a7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10815, 'h10825, 'h109a8, 'h10835, 'h10845, 'h109a9, 'h10ba5, 'h10855, 'h10865, 'h109aa, 'h10875, 'h10885, 'h109ab, 'h10895, 'h103bc, 'h108a5, 'h109ac, 'h108b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c5, 'h109ad, 'h108d5, 'h106e5, 'h109ae, 'h10bb5, 'h106f5, 'h10705, 'h109af, 'h10715, 'h10725, 'h109b0, 'h10735, 'h10745, 'h109b1, 'h103bc, 'h10755, 'h10765, 'h109b2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10775, 'h10785, 'h109b3, 'h10795, 'h10bb5, 'h107a5, 'h109b4, 'h107b5, 'h107c5, 'h109b5, 'h107d5, 'h107e5, 'h109b6, 'h107f5, 'h103bc, 'h10805, 'h109b7, 'h10815, 'h21f8e, 'h21f8f, 'h21f8d, 'h10825, 'h109b8, 'h10835, 'h10845, 'h109b9, 'h10bb5, 'h10855, 'h10865, 'h109ba, 'h10875, 'h10885, 'h109bb, 'h10895, 'h108a5, 'h109bc, 'h103bc, 'h108b5, 'h108c5, 'h109bd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d5, 'h106e5, 'h109be, 'h10bc5, 'h106f5, 'h10705, 'h109bf, 'h10715, 'h10725, 'h109c0, 'h10735, 'h10745, 'h109c1, 'h10755, 'h103bc, 'h10765, 'h109c2, 'h10775, 'h21f8e, 'h21f8f, 'h21f8d, 'h10785, 'h109c3, 'h10795, 'h10bc5, 'h107a5, 'h109c4, 'h107b5, 'h107c5, 'h109c5, 'h107d5, 'h107e5, 'h109c6, 'h107f5, 'h10805, 'h109c7, 'h103bc, 'h10815, 'h10825, 'h109c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10835, 'h10845, 'h109c9, 'h10bc5, 'h10855, 'h10865, 'h109ca, 'h10875, 'h10885, 'h109cb, 'h10895, 'h108a5, 'h109cc, 'h108b5, 'h103bc, 'h108c5, 'h109cd, 'h108d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h109ce, 'h10bd5, 'h106f5, 'h10705, 'h109cf, 'h10715, 'h10725, 'h109d0, 'h10735, 'h10745, 'h109d1, 'h10755, 'h10765, 'h109d2, 'h103bc};
	int DATA4 [4*SIZE-1:0] = {DATA3, DATA0};
	
endpackage
