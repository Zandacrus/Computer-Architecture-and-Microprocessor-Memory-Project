

package LU_PKG_2;
	
	import LU_PKG_1::DATA1;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h100154, 'h100155, 'h1000d0, 'h100156, 'h1000d1, 'h100157, 'h1000d2, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h10003c, 'h2004f7, 'h100160, 'h1000d3, 'h100047, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h1000d0, 'h100166, 'h1000d1, 'h100167, 'h1000d2, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10003c, 'h2004f7, 'h10016e, 'h10016f, 'h100047, 'h100170, 'h1000d3, 'h1000d8, 'h1000d7, 'h1000d4, 'h1000d9, 'h1000d5, 'h1000da, 'h1000d6, 'h1000db, 'h1000dc, 'h1000dd, 'h1000de, 'h1000df, 'h1000e0, 'h1000e1, 'h10003c, 'h2004f7, 'h1000e2, 'h1000e3, 'h100047, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000d7, 'h1000e8, 'h1000d4, 'h1000e9, 'h1000d5, 'h1000ea, 'h1000d6, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h10003c, 'h2004f7, 'h1000f0, 'h1000f1, 'h100047, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000d7, 'h1000f8, 'h1000d4, 'h1000f9, 'h1000d5, 'h1000fa, 'h1000d6, 'h1000fb, 'h1000fc, 'h1000fd, 'h10003c, 'h2004f7, 'h1000fe, 'h1000ff, 'h100047, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h1000d7, 'h100108, 'h1000d4, 'h100109, 'h1000d5, 'h10010a, 'h1000d6, 'h10010b, 'h10003c, 'h2004f7, 'h10010c, 'h10010d, 'h100047, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h1000d7, 'h100118, 'h1000d4, 'h100119, 'h1000d5, 'h10011a, 'h10003c, 'h2004f7, 'h1000d6, 'h10011b, 'h100047, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h1000d7, 'h100128, 'h1000d4, 'h100129, 'h10003c, 'h2004f7, 'h1000d5, 'h10012a, 'h100047, 'h1000d6, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h1000d7, 'h100138, 'h10003c, 'h2004f7, 'h1000d4, 'h100139, 'h100047, 'h1000d5, 'h10013a, 'h1000d6, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h1000d7, 'h100146, 'h10003c, 'h2004f7, 'h100147, 'h100148, 'h100047, 'h100149, 'h1000d4, 'h1000d5, 'h10014a, 'h1000d6, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h1000d7, 'h100154, 'h10003c, 'h2004f7, 'h100155, 'h100156, 'h100047, 'h100157, 'h100158, 'h100159, 'h1000d4, 'h10015a, 'h1000d5, 'h10015b, 'h1000d6, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h1000d7, 'h100162, 'h10003c, 'h2004f7, 'h100163, 'h100164, 'h100047, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h1000d4, 'h10016a, 'h1000d5, 'h10016b, 'h1000d6, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h1000d7, 'h10003c, 'h2004f7, 'h1000dc, 'h1000db, 'h100047, 'h1000d8, 'h1000dd, 'h1000d9, 'h1000de, 'h1000da, 'h1000df, 'h1000e0, 'h1000e1, 'h1000e2, 'h1000e3, 'h1000e4, 'h1000e5, 'h1000e6, 'h1000e7, 'h1000e8, 'h1000e9, 'h10003c, 'h2004f7, 'h1000ea, 'h1000eb, 'h100047, 'h1000db, 'h1000ec, 'h1000d8, 'h1000ed, 'h1000d9, 'h1000ee, 'h1000da, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h10003c, 'h2004f7, 'h1000f8, 'h1000f9, 'h100047, 'h1000fa, 'h1000fb, 'h1000db, 'h1000fc, 'h1000d8, 'h1000fd, 'h1000d9, 'h1000fe, 'h1000da, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100105, 'h10003c, 'h2004f7, 'h100106, 'h100107, 'h100047, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h1000db, 'h10010c, 'h1000d8, 'h10010d, 'h1000d9, 'h10010e, 'h1000da, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h10003c, 'h2004f7, 'h100114, 'h100115, 'h100047, 'h100116, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h1000db, 'h10011c, 'h1000d8, 'h10011d, 'h1000d9, 'h10011e, 'h1000da, 'h10011f, 'h100120, 'h100121, 'h10003c, 'h2004f7, 'h100122, 'h100123, 'h100047, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h1000db, 'h10012c, 'h1000d8, 'h10012d, 'h1000d9, 'h10012e, 'h1000da, 'h10012f, 'h10003c, 'h2004f7, 'h100130, 'h100131, 'h100047, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h1000db, 'h10013c, 'h10013d, 'h1000d8, 'h1000d9, 'h10013e, 'h10003c, 'h2004f7, 'h1000da, 'h10013f, 'h100047, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h1000db, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h1000d8, 'h10003c, 'h2004f7, 'h1000d9, 'h10014e, 'h100047, 'h1000da, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h1000db, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10003c, 'h2004f7, 'h10015d, 'h1000d8, 'h100047, 'h10015e, 'h1000d9, 'h10015f, 'h1000da, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h1000db, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10003c, 'h2004f7, 'h10016b, 'h10016c, 'h100047, 'h10016d, 'h1000d8, 'h10016e, 'h1000d9, 'h10016f, 'h1000da, 'h100170, 'h1000e0, 'h1000df, 'h1000e1, 'h1000dc, 'h1000dd, 'h1000e2, 'h1000de, 'h1000e3, 'h1000e4, 'h1000e5, 'h10003c, 'h2004f7, 'h1000e6, 'h100047, 'h1000e7, 'h1000e8, 'h1000e9, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h1000df, 'h1000f0, 'h1000f1, 'h1000dc, 'h1000dd, 'h1000f2, 'h1000de, 'h1000f3, 'h10003c, 'h2004f7, 'h1000f4, 'h1000f5, 'h100047, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000df, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h1000dc, 'h1000dd, 'h100102, 'h10003c, 'h2004f7, 'h1000de, 'h100103, 'h100047, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h1000df, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h1000dc, 'h10003c, 'h2004f7, 'h1000dd, 'h100112, 'h100047, 'h1000de, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h100119, 'h1000df, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h10003c, 'h2004f7, 'h1000dc, 'h100047, 'h1000dd, 'h100122, 'h1000de, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h1000df, 'h100128, 'h10012a, 'h100129, 'h10012b, 'h10012c, 'h10012e, 'h10012d, 'h10012f, 'h10003c, 'h2004f7, 'h100130, 'h100047, 'h100132, 'h1000dc, 'h100131, 'h1000dd, 'h1000de, 'h100133, 'h100134, 'h100136, 'h1000df, 'h100135, 'h100137, 'h100138, 'h10013a, 'h100139, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10003c, 'h2004f7, 'h100047, 'h10013f, 'h100140, 'h100141, 'h100142, 'h1000dc, 'h1000dd, 'h1000de, 'h100143, 'h1000df, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10003c, 'h2004f7, 'h100047, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h1000dc, 'h1000dd, 'h1000de, 'h100153, 'h1000df, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10003c, 'h2004f7, 'h100047, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h1000dc, 'h1000dd, 'h100163, 'h1000de, 'h100164, 'h1000df, 'h100165, 'h100166, 'h100167, 'h100168, 'h10003c, 'h2004f7, 'h100047, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h1000e4, 'h1000e3, 'h1000e0, 'h1000e5, 'h1000e1, 'h1000e6, 'h1000e2, 'h1000e7, 'h1000e8, 'h1000e9, 'h10003c, 'h2004f7, 'h100047, 'h1000ea, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000e3, 'h1000f4, 'h1000e0, 'h1000f5, 'h1000e1, 'h1000f6, 'h1000e2, 'h1000f7, 'h10003c, 'h2004f7, 'h100047, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h1000e3, 'h100104, 'h1000e0, 'h100105, 'h1000e1, 'h100106, 'h10003c, 'h2004f7, 'h100047, 'h1000e2, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h1000e3, 'h100114, 'h1000e0, 'h100115, 'h10003c, 'h2004f7, 'h100047, 'h1000e1, 'h100116, 'h1000e2, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h1000e3, 'h100124, 'h10003c, 'h2004f7, 'h100047, 'h1000e0, 'h100125, 'h1000e1, 'h100126, 'h1000e2, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h10003c, 'h2004f7, 'h100047, 'h1000e3, 'h100134, 'h100135, 'h1000e0, 'h1000e1, 'h100136, 'h1000e2, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h10003c, 'h2004f7, 'h100047, 'h1000e3, 'h100142, 'h100143, 'h100144, 'h100145, 'h1000e0, 'h1000e1, 'h100146, 'h1000e2, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h10003c, 'h2004f7, 'h100047, 'h1000e3, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h1000e0, 'h1000e1, 'h100156, 'h1000e2, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10003c, 'h2004f7, 'h100047, 'h1000e3, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h1000e0, 'h100166, 'h1000e1, 'h100167, 'h1000e2, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10003c, 'h2004f7, 'h100047, 'h10016c, 'h1000e3, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h1000e8, 'h1000e7, 'h1000e4, 'h1000e9, 'h1000e5, 'h1000ea, 'h1000e6, 'h1000eb, 'h1000ec, 'h1000ed, 'h1000ee, 'h1000ef, 'h10003c, 'h2004f7, 'h100047, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000e7, 'h1000f8, 'h1000e4, 'h1000f9, 'h1000e5, 'h1000fa, 'h1000e6, 'h1000fb, 'h1000fc, 'h1000fd, 'h10003c, 'h2004f7, 'h100047, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h1000e7, 'h100108, 'h1000e4, 'h100109, 'h1000e5, 'h10010a, 'h1000e6, 'h10010b, 'h10003c, 'h2004f7, 'h100047, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h1000e7, 'h100118, 'h1000e4, 'h100119, 'h1000e5, 'h10011a, 'h10003c, 'h2004f7, 'h100047, 'h1000e6, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h1000e7, 'h100128, 'h1000e4, 'h100129, 'h10003c, 'h2004f7, 'h100047, 'h1000e5, 'h10012a, 'h1000e6, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h1000e7, 'h100136, 'h100137, 'h100138, 'h10003c, 'h2004f7, 'h100047, 'h100139, 'h1000e4, 'h1000e5, 'h10013a, 'h1000e6, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h1000e7, 'h100144, 'h100145, 'h100146, 'h10003c, 'h2004f7, 'h100047, 'h100147, 'h100148, 'h100149, 'h1000e4, 'h1000e5, 'h10014a, 'h1000e6, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h1000e7, 'h100152, 'h100153, 'h100154, 'h10003c, 'h2004f7, 'h100047, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h1000e4, 'h1000e5, 'h10015a, 'h1000e6, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h1000e7, 'h100160, 'h100161, 'h100162, 'h10003c, 'h2004f7, 'h100047, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h1000e4, 'h10016a, 'h1000e5, 'h10016b, 'h1000e6, 'h10016c, 'h10016d, 'h1000e7, 'h10016e, 'h10016f, 'h100170, 'h10003c, 'h2004f7, 'h100047, 'h1000ec, 'h1000eb, 'h1000e8, 'h1000ed, 'h1000e9, 'h1000ee, 'h1000ea, 'h1000ef, 'h1000f0, 'h1000f1, 'h1000f2, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h1000f7, 'h1000f8, 'h1000f9, 'h10003c, 'h2004f7, 'h100047, 'h1000fa, 'h1000fb, 'h1000eb, 'h1000fc, 'h1000e8, 'h1000fd, 'h1000e9, 'h1000fe, 'h1000ea, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h10003c, 'h2004f7, 'h100047, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h1000eb, 'h10010c, 'h1000e8, 'h10010d, 'h1000e9, 'h10010e, 'h1000ea, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100114, 'h100115, 'h10003c, 'h2004f7, 'h100047, 'h100116, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h1000eb, 'h10011c, 'h1000e8, 'h10011d, 'h1000e9, 'h10011e, 'h1000ea, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h10003c, 'h2004f7, 'h100047, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h1000eb, 'h10012c, 'h10012d, 'h1000e8, 'h1000e9, 'h10012e, 'h1000ea, 'h10012f, 'h100130, 'h100131, 'h10003c, 'h2004f7, 'h100047, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h1000eb, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h1000e8, 'h1000e9, 'h10013e, 'h1000ea, 'h10013f, 'h10003c, 'h2004f7, 'h100047, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h1000eb, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h1000e8, 'h1000e9, 'h10014e, 'h10003c, 'h2004f7, 'h100047, 'h1000ea, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h1000eb, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h1000e8, 'h10003c, 'h2004f7, 'h100047, 'h1000e9, 'h10015e, 'h1000ea, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h1000eb, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10003c, 'h2004f7, 'h100047, 'h10016d, 'h1000e8, 'h10016e, 'h1000e9, 'h10016f, 'h1000ea, 'h100170, 'h1000f0, 'h1000ef, 'h1000ec, 'h1000f1, 'h1000ed, 'h1000f2, 'h1000ee, 'h1000f3, 'h1000f4, 'h1000f5, 'h1000f6, 'h10003c, 'h2004f7, 'h100047, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h1000ef, 'h100100, 'h1000ec, 'h100101, 'h1000ed, 'h100102, 'h1000ee, 'h100103, 'h100104, 'h10003c, 'h2004f7, 'h100047, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h1000ef, 'h100110, 'h1000ec, 'h100111, 'h1000ed, 'h100112, 'h1000ee, 'h10003c, 'h2004f7, 'h100047, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h1000ef, 'h100120, 'h1000ec, 'h100121, 'h1000ed, 'h10003c, 'h2004f7, 'h100047, 'h100122, 'h1000ee, 'h100123, 'h100124, 'h100125, 'h100126, 'h100127, 'h100128, 'h100129, 'h10012a, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h1000ef, 'h100130, 'h100131, 'h1000ec, 'h10003c, 'h2004f7, 'h100047, 'h1000ed, 'h100132, 'h1000ee, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h1000ef, 'h10013e, 'h10013f, 'h100140, 'h10003c, 'h2004f7, 'h100047, 'h100141, 'h1000ec, 'h1000ed, 'h100142, 'h1000ee, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h1000ef, 'h10014c, 'h10014d, 'h10014e, 'h10003c, 'h2004f7, 'h100047, 'h10014f, 'h100150, 'h100151, 'h1000ec, 'h1000ed, 'h100152, 'h1000ee, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h1000ef, 'h10015a, 'h10015b, 'h10015c, 'h10003c, 'h2004f7, 'h100047, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h1000ec, 'h1000ed, 'h100162, 'h1000ee, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h1000ef, 'h100168, 'h100169, 'h10016a, 'h10003c, 'h2004f7, 'h100047, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h1000f4, 'h1000f3, 'h1000f0, 'h1000f5, 'h1000f1, 'h1000f6, 'h1000f2, 'h1000f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1000fb, 'h10003c, 'h2004f7, 'h100047, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h1000f3, 'h100104, 'h1000f0, 'h100105, 'h1000f1, 'h100106, 'h1000f2, 'h100107, 'h100108, 'h100109, 'h10003c, 'h2004f7, 'h100047, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h1000f3, 'h100114, 'h1000f0, 'h100115, 'h1000f1, 'h100116, 'h1000f2, 'h100117, 'h10003c, 'h2004f7, 'h100047, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h100122, 'h100123, 'h1000f3, 'h100124, 'h100125, 'h1000f0, 'h1000f1, 'h100126, 'h10003c, 'h2004f7, 'h100047, 'h1000f2, 'h100127, 'h100129, 'h10012a, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h1000f3, 'h100134, 'h100135, 'h1000f0, 'h1000f1, 'h100136, 'h10003c, 'h2004f7, 'h100047, 'h1000f2, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h1000f3, 'h100142, 'h100143, 'h100144, 'h100145, 'h1000f0, 'h10003c, 'h2004f7, 'h100047, 'h1000f1, 'h100146, 'h1000f2, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h1000f3, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h10003c, 'h2004f7, 'h100047, 'h100155, 'h1000f0, 'h1000f1, 'h100156, 'h1000f2, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h1000f3, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h10003c, 'h2004f7, 'h100047, 'h100163, 'h100164, 'h100165, 'h1000f0, 'h1000f1, 'h100166, 'h1000f2, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h1000f3, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h10003c, 'h2004f7, 'h100047, 'h1000f8, 'h1000f7, 'h1000f4, 'h1000f9, 'h1000f5, 'h1000fa, 'h1000f6, 'h1000fb, 'h1000fc, 'h1000fd, 'h1000fe, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h100103, 'h100104, 'h100105, 'h10003c, 'h2004f7, 'h100047, 'h100106, 'h100107, 'h1000f7, 'h100108, 'h1000f4, 'h100109, 'h1000f5, 'h10010a, 'h1000f6, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h10003c, 'h2004f7, 'h100047, 'h100114, 'h100115, 'h100116, 'h100117, 'h1000f7, 'h100118, 'h1000f4, 'h100119, 'h1000f5, 'h10011a, 'h1000f6, 'h10011b, 'h10011c, 'h10011d, 'h10011e, 'h10011f, 'h100120, 'h100121, 'h10003c, 'h2004f7, 'h100047, 'h100122, 'h100123, 'h100125, 'h100126, 'h100127, 'h1000f7, 'h100129, 'h1000f4, 'h1000f5, 'h10012a, 'h1000f6, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h10003c, 'h2004f7, 'h100047, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h1000f7, 'h100138, 'h100139, 'h1000f4, 'h1000f5, 'h10013a, 'h1000f6, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h10003c, 'h2004f7, 'h100047, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h1000f7, 'h100146, 'h100147, 'h100148, 'h100149, 'h1000f4, 'h1000f5, 'h10014a, 'h1000f6, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10003c, 'h2004f7, 'h100047, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h1000f7, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h1000f4, 'h1000f5, 'h10015a, 'h1000f6, 'h10015b, 'h10015c, 'h10003c, 'h2004f7, 'h100047, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h1000f7, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h1000f4, 'h1000f5, 'h10016a, 'h1000f6, 'h10003c, 'h2004f7, 'h100047, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h1000f7, 'h100170, 'h1000fc, 'h1000fb, 'h1000fd, 'h1000f8, 'h1000f9, 'h1000fe, 'h1000fa, 'h1000ff, 'h100100, 'h100101, 'h100102, 'h10003c, 'h2004f7, 'h100047, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h1000fb, 'h10010c, 'h10010d, 'h1000f8, 'h1000f9, 'h10010e, 'h1000fa, 'h10010f, 'h100110, 'h100112, 'h10003c, 'h2004f7, 'h100047, 'h100111, 'h100113, 'h100114, 'h100116, 'h100115, 'h100117, 'h100118, 'h10011a, 'h1000fb, 'h100119, 'h10011b, 'h10011c, 'h10011e, 'h10011d, 'h1000f8, 'h1000f9, 'h1000fa, 'h10011f, 'h10003c, 'h2004f7, 'h100047, 'h100121, 'h100122, 'h100123, 'h100125, 'h100126, 'h100127, 'h100129, 'h10012a, 'h1000fb, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h1000f8, 'h1000f9, 'h10003c, 'h2004f7, 'h100047, 'h1000fa, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h1000fb, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h10003c, 'h2004f7, 'h100047, 'h1000f8, 'h1000f9, 'h1000fa, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h1000fb, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h10003c, 'h2004f7, 'h100047, 'h100151, 'h100152, 'h1000f8, 'h1000f9, 'h1000fa, 'h100153, 'h100154, 'h100155, 'h1000fb, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10003c, 'h2004f7, 'h100047, 'h10015f, 'h100160, 'h100161, 'h100162, 'h1000f8, 'h1000f9, 'h1000fa, 'h100163, 'h1000fb, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10003c, 'h2004f7, 'h100047, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h100100, 'h1000ff, 'h1000fc, 'h100101, 'h1000fd, 'h100102, 'h1000fe, 'h100103, 'h100104, 'h100105, 'h100106, 'h100107, 'h100108, 'h100109, 'h10003c, 'h2004f7, 'h100047, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h1000ff, 'h100110, 'h1000fc, 'h100111, 'h1000fd, 'h100112, 'h1000fe, 'h100113, 'h100114, 'h100115, 'h100116, 'h100117, 'h10003c, 'h2004f7, 'h100047, 'h100118, 'h100119, 'h10011a, 'h10011b, 'h10011d, 'h10011e, 'h10011f, 'h1000ff, 'h100121, 'h1000fc, 'h1000fd, 'h100122, 'h1000fe, 'h100123, 'h100125, 'h100126, 'h100127, 'h100129, 'h10003c, 'h2004f7, 'h100047, 'h10012a, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h1000ff, 'h100132, 'h100133, 'h100134, 'h100135, 'h1000fc, 'h1000fd, 'h100136, 'h1000fe, 'h100137, 'h100138, 'h10003c, 'h2004f7, 'h100047, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h1000ff, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h1000fc, 'h1000fd, 'h100146, 'h1000fe, 'h10003c, 'h2004f7, 'h100047, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h1000ff, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h1000fc, 'h1000fd, 'h10003c, 'h2004f7, 'h100047, 'h100156, 'h1000fe, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h1000ff, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h10003c, 'h2004f7, 'h100047, 'h1000fc, 'h1000fd, 'h100166, 'h1000fe, 'h100167, 'h100168, 'h100169, 'h1000ff, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h100104, 'h100103, 'h100100, 'h10003c, 'h2004f7, 'h100047, 'h100105, 'h100101, 'h100106, 'h100102, 'h100107, 'h100108, 'h100109, 'h10010a, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h100113, 'h100103, 'h10003c, 'h2004f7, 'h100047, 'h100114, 'h100115, 'h100100, 'h100101, 'h100116, 'h100102, 'h100117, 'h100119, 'h10011a, 'h10011b, 'h10011d, 'h10011e, 'h10011f, 'h100121, 'h100122, 'h100123, 'h100125, 'h100103, 'h10003c, 'h2004f7, 'h100047, 'h100126, 'h100127, 'h100129, 'h100100, 'h100101, 'h10012a, 'h100102, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100103, 'h10003c, 'h2004f7, 'h100047, 'h100136, 'h100137, 'h100138, 'h100139, 'h100100, 'h100101, 'h10013a, 'h100102, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100103, 'h10003c, 'h2004f7, 'h100047, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h100100, 'h100101, 'h10014a, 'h100102, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100103, 'h10003c, 'h2004f7, 'h100047, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h100100, 'h100101, 'h10015a, 'h100102, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100103, 'h10003c, 'h2004f7, 'h100047, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h100100, 'h100101, 'h10016a, 'h100102, 'h10016b, 'h10016c, 'h10016d, 'h100103, 'h10003c, 'h2004f7, 'h100047, 'h10016e, 'h10016f, 'h100170, 'h100108, 'h100107, 'h100104, 'h100109, 'h100105, 'h10010a, 'h100106, 'h10010b, 'h10010c, 'h10010d, 'h10010e, 'h10010f, 'h100110, 'h100111, 'h100112, 'h10003c, 'h2004f7, 'h100047, 'h100113, 'h100115, 'h100116, 'h100117, 'h100107, 'h100119, 'h100104, 'h100105, 'h10011a, 'h100106, 'h10011b, 'h10011d, 'h10011e, 'h10011f, 'h100121, 'h100122, 'h100123, 'h100125, 'h10003c, 'h2004f7, 'h100047, 'h100126, 'h100127, 'h100129, 'h10012a, 'h10012b, 'h100107, 'h10012d, 'h100104, 'h100105, 'h10012e, 'h100106, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h10003c, 'h2004f7, 'h100047, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h100107, 'h10013c, 'h10013d, 'h100104, 'h100105, 'h10013e, 'h100106, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h10003c, 'h2004f7, 'h100047, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h100107, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h100104, 'h100105, 'h10014e, 'h100106, 'h10014f, 'h100150, 'h100151, 'h10003c, 'h2004f7, 'h100047, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100107, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h100104, 'h100105, 'h10015e, 'h100106, 'h10015f, 'h10003c, 'h2004f7, 'h100047, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100107, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h100104, 'h100105, 'h10016e, 'h10003c, 'h2004f7, 'h100047, 'h100106, 'h10016f, 'h100170, 'h10010c, 'h10010b, 'h10010d, 'h100108, 'h100109, 'h10010e, 'h10010a, 'h10010f, 'h100111, 'h100112, 'h100113, 'h100115, 'h100116, 'h100117, 'h100119, 'h10003c, 'h2004f7, 'h100047, 'h10011a, 'h10011b, 'h10011d, 'h10011e, 'h10011f, 'h10010b, 'h100121, 'h100108, 'h100109, 'h100122, 'h10010a, 'h100123, 'h100125, 'h100126, 'h100127, 'h100129, 'h10012a, 'h10012b, 'h10003c, 'h2004f7, 'h100047, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h10010b, 'h100132, 'h100133, 'h100134, 'h100135, 'h100108, 'h100109, 'h100136, 'h10010a, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10003c, 'h2004f7, 'h100047, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h10010b, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100108, 'h100109, 'h100146, 'h10010a, 'h100147, 'h100148, 'h10003c, 'h2004f7, 'h100047, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10010b, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100108, 'h100109, 'h100156, 'h10010a, 'h10003c, 'h2004f7, 'h100047, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10010b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100108, 'h100109, 'h10003c, 'h2004f7, 'h100047, 'h100166, 'h10010a, 'h100167, 'h100168, 'h100169, 'h10010b, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h100111, 'h10010f, 'h10010d, 'h100112, 'h10010e, 'h10003c, 'h2004f7, 'h100047, 'h100113, 'h100115, 'h100116, 'h100117, 'h100119, 'h10011a, 'h10011b, 'h10011d, 'h10011e, 'h10011f, 'h100121, 'h100122, 'h100123, 'h100125, 'h10010f, 'h10010d, 'h100126, 'h10010e, 'h10003c, 'h2004f7, 'h100047, 'h100127, 'h100129, 'h10012a, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h10010f, 'h100138, 'h100139, 'h10003c, 'h2004f7, 'h100047, 'h10010d, 'h10013a, 'h10010e, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h10010f, 'h100148, 'h10003c, 'h2004f7, 'h100047, 'h100149, 'h10010d, 'h10014a, 'h10010e, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h10010f, 'h10003c, 'h2004f7, 'h100047, 'h100158, 'h100159, 'h10010d, 'h10015a, 'h10010e, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h10003c, 'h2004f7, 'h100047, 'h10010f, 'h100168, 'h100169, 'h10010d, 'h10016a, 'h10010e, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h100115, 'h100113, 'h100111, 'h100116, 'h100112, 'h100117, 'h10003c, 'h2004f7, 'h100047, 'h100119, 'h10011a, 'h10011b, 'h10011d, 'h10011e, 'h10011f, 'h100121, 'h100122, 'h100123, 'h100125, 'h100126, 'h100127, 'h100129, 'h100113, 'h100111, 'h10012a, 'h100112, 'h10012b, 'h10003c, 'h2004f7, 'h100047, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h100113, 'h100111, 'h10013a, 'h100112, 'h10013b, 'h10003c, 'h2004f7, 'h100047, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100113, 'h100149, 'h100111, 'h10014a, 'h100112, 'h10003c, 'h2004f7, 'h100047, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100113, 'h100158, 'h100159, 'h100111, 'h10015a, 'h10003c, 'h2004f7, 'h100047, 'h100112, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100113, 'h100168, 'h100169, 'h100111, 'h10003c, 'h2004f7, 'h100047, 'h10016a, 'h100112, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h100119, 'h100117, 'h100115, 'h10011a, 'h100116, 'h10011b, 'h10011d, 'h10011e, 'h10011f, 'h100121, 'h10003c, 'h2004f7, 'h100047, 'h100122, 'h100123, 'h100125, 'h100126, 'h100127, 'h100129, 'h10012a, 'h10012b, 'h10012d, 'h100117, 'h100115, 'h10012e, 'h100116, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h10003c, 'h2004f7, 'h100047, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h100117, 'h10013d, 'h100115, 'h10013e, 'h100116, 'h10013f, 'h100140, 'h100141, 'h100142, 'h10003c, 'h2004f7, 'h100047, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h100117, 'h10014c, 'h10014d, 'h100115, 'h10014e, 'h100116, 'h10014f, 'h100150, 'h100151, 'h10003c, 'h2004f7, 'h100047, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h100117, 'h10015c, 'h10015d, 'h100115, 'h10015e, 'h100116, 'h10015f, 'h100160, 'h10003c, 'h2004f7, 'h100047, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h100117, 'h10016c, 'h10016d, 'h100115, 'h10016e, 'h100116, 'h10016f, 'h10003c, 'h2004f7, 'h100047, 'h100170, 'h10011d, 'h10011b, 'h100119, 'h10011e, 'h10011a, 'h10011f, 'h100121, 'h100122, 'h100123, 'h100125, 'h100126, 'h100127, 'h100129, 'h10012a, 'h10012b, 'h10012d, 'h10012e, 'h10003c, 'h2004f7, 'h100047, 'h10012f, 'h100130, 'h10011b, 'h100131, 'h100119, 'h100132, 'h10011a, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10003c, 'h2004f7, 'h100047, 'h10013e, 'h10013f, 'h10011b, 'h100140, 'h100141, 'h100119, 'h100142, 'h10011a, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10003c, 'h2004f7, 'h100047, 'h10014d, 'h10014e, 'h10014f, 'h10011b, 'h100150, 'h100151, 'h100119, 'h100152, 'h10011a, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10003c, 'h2004f7, 'h100047, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h10011b, 'h100160, 'h100161, 'h100119, 'h100162, 'h10011a, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10003c, 'h2004f7, 'h100047, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h10011b, 'h100170, 'h100121, 'h10011f, 'h10011d, 'h100122, 'h10011e, 'h100123, 'h100125, 'h100126, 'h100127, 'h100129, 'h10012a, 'h10003c, 'h2004f7, 'h100047, 'h10012b, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h100131, 'h100132, 'h100133, 'h10011f, 'h100134, 'h100135, 'h10011d, 'h100136, 'h10011e, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10003c, 'h2004f7, 'h100047, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h10011f, 'h100144, 'h100145, 'h10011d, 'h100146, 'h10011e, 'h100147, 'h100148, 'h100149, 'h10003c, 'h2004f7, 'h100047, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h10011f, 'h100154, 'h100155, 'h10011d, 'h100156, 'h10011e, 'h100157, 'h100158, 'h10003c, 'h2004f7, 'h100047, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h10011f, 'h100164, 'h100165, 'h10011d, 'h100166, 'h10011e, 'h100167, 'h10003c, 'h2004f7, 'h100047, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h100125, 'h100123, 'h100127, 'h100121, 'h100126, 'h100122, 'h100129, 'h10012b, 'h10012a, 'h10003c, 'h2004f7, 'h100047, 'h10012d, 'h10012f, 'h10012e, 'h100130, 'h100131, 'h100133, 'h100132, 'h100134, 'h100135, 'h100137, 'h100123, 'h100136, 'h100121, 'h100138, 'h100139, 'h10013b, 'h10013a, 'h100122, 'h10003c, 'h2004f7, 'h100047, 'h10013c, 'h10013d, 'h10013f, 'h10013e, 'h100140, 'h100141, 'h100143, 'h100142, 'h100144, 'h100145, 'h100123, 'h100147, 'h100121, 'h100146, 'h100148, 'h100149, 'h10014b, 'h10014a, 'h10003c, 'h2004f7, 'h100047, 'h100122, 'h10014c, 'h10014d, 'h10014f, 'h10014e, 'h100150, 'h100151, 'h100153, 'h100152, 'h100154, 'h100123, 'h100155, 'h100157, 'h100121, 'h100156, 'h100158, 'h100159, 'h10015b, 'h10003c, 'h2004f7, 'h100047, 'h10015a, 'h100122, 'h10015c, 'h10015d, 'h10015f, 'h10015e, 'h100160, 'h100161, 'h100163, 'h100162, 'h100123, 'h100164, 'h100165, 'h100167, 'h100121, 'h100166, 'h100168, 'h100169, 'h10016b, 'h10003c, 'h2004f7, 'h100047, 'h10016a, 'h100122, 'h10016c, 'h10016d, 'h10016f, 'h10016e, 'h100170, 'h100129, 'h100127, 'h100125, 'h10012a, 'h100126, 'h10012b, 'h10012c, 'h10012d, 'h10012e, 'h10012f, 'h100130, 'h10003c, 'h2004f7, 'h100047, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100127, 'h100139, 'h100125, 'h10013a, 'h100126, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h10003c, 'h2004f7, 'h100047, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100127, 'h100148, 'h100149, 'h100125, 'h10014a, 'h100126, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10003c, 'h2004f7, 'h100047, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100127, 'h100158, 'h100159, 'h100125, 'h10015a, 'h100126, 'h10015b, 'h10015c, 'h10015d, 'h10003c, 'h2004f7, 'h100047, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100127, 'h100168, 'h100169, 'h100125, 'h10016a, 'h100126, 'h10016b, 'h10016c, 'h10003c, 'h2004f7, 'h100047, 'h10016d, 'h10016e, 'h10016f, 'h100170, 'h10012d, 'h10012c, 'h100129, 'h10012e, 'h10012a, 'h10012f, 'h10012b, 'h100130, 'h100131, 'h100132, 'h100133, 'h100134, 'h100135, 'h100136, 'h10003c, 'h2004f7, 'h100047, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10012c, 'h100129, 'h10013e, 'h10012a, 'h10013f, 'h10012b, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h10003c, 'h2004f7, 'h100047, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10012c, 'h100129, 'h10014e, 'h10012a, 'h10014f, 'h10012b, 'h100150, 'h100151, 'h100152, 'h10003c, 'h2004f7, 'h100047, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10012c, 'h100129, 'h10015e, 'h10012a, 'h10015f, 'h10012b, 'h100160, 'h10003c, 'h2004f7, 'h100047, 'h100161, 'h100162, 'h100163, 'h100164, 'h100165, 'h100166, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016d, 'h10012c, 'h10016e, 'h100129, 'h10012a, 'h10016f, 'h10003c, 'h2004f7, 'h100047, 'h10012b, 'h100170, 'h100131, 'h100130, 'h10012d, 'h100132, 'h10012e, 'h100133, 'h10012f, 'h100134, 'h100135, 'h100136, 'h100137, 'h100138, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10003c, 'h2004f7, 'h100047, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100130, 'h100141, 'h10012d, 'h100142, 'h10012e, 'h100143, 'h10012f, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10003c, 'h2004f7, 'h100047, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100130, 'h100151, 'h10012d, 'h100152, 'h10012e, 'h100153, 'h10012f, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h10003c, 'h2004f7, 'h100047, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100130, 'h100161, 'h10012d, 'h100162, 'h10012e, 'h100163, 'h10012f, 'h100164, 'h100165, 'h100166, 'h10003c, 'h2004f7, 'h100047, 'h100167, 'h100168, 'h100169, 'h10016a, 'h10016b, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h100130, 'h100135, 'h100134, 'h100131, 'h100136, 'h100132, 'h100137, 'h100133, 'h100138, 'h10003c, 'h2004f7, 'h100047, 'h100139, 'h10013a, 'h10013b, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100134, 'h100145, 'h100131, 'h100146, 'h100132, 'h100147, 'h10003c, 'h2004f7, 'h100047, 'h100133, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100134, 'h100155, 'h100131, 'h100156, 'h10003c, 'h2004f7, 'h100047, 'h100132, 'h100157, 'h100133, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100134, 'h100165, 'h10003c, 'h2004f7, 'h100047, 'h100166, 'h100131, 'h100132, 'h100167, 'h100133, 'h100168, 'h10016a, 'h10016b, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h100139, 'h100138, 'h100135, 'h10013a, 'h100136, 'h10013b, 'h10003c, 'h2004f7, 'h100047, 'h100137, 'h10013c, 'h10013d, 'h10013e, 'h10013f, 'h100140, 'h100141, 'h100142, 'h100143, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100138, 'h100149, 'h100135, 'h10014a, 'h10003c, 'h2004f7, 'h100047, 'h100136, 'h10014b, 'h100137, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100138, 'h100159, 'h10003c, 'h2004f7, 'h100047, 'h100135, 'h10015a, 'h100136, 'h10015b, 'h100137, 'h10015c, 'h10015d, 'h10015e, 'h10015f, 'h100160, 'h100161, 'h100162, 'h100163, 'h100164, 'h100166, 'h100167, 'h100168, 'h100138, 'h10003c, 'h2004f7, 'h100047, 'h10016a, 'h100135, 'h100136, 'h10016b, 'h100137, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h10013d, 'h10013c, 'h10013f, 'h100139, 'h10013e, 'h10013a, 'h10013b, 'h100140, 'h100141, 'h100143, 'h10003c, 'h2004f7, 'h100047, 'h100142, 'h100144, 'h100145, 'h100147, 'h100146, 'h100148, 'h100149, 'h10014b, 'h10014a, 'h10014c, 'h10013c, 'h10014d, 'h10014f, 'h100139, 'h10014e, 'h10013a, 'h10013b, 'h100150, 'h10003c, 'h2004f7, 'h100047, 'h100151, 'h100153, 'h100152, 'h100154, 'h100155, 'h100157, 'h100156, 'h100158, 'h100159, 'h10015b, 'h10013c, 'h10015a, 'h10015c, 'h10015d, 'h10015f, 'h10015e, 'h100139, 'h10013a, 'h10003c, 'h2004f7, 'h100047, 'h10013b, 'h100160, 'h100162, 'h100163, 'h100164, 'h100166, 'h100167, 'h100168, 'h10016a, 'h10016b, 'h10013c, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h100141, 'h100140, 'h10013d, 'h10003c, 'h2004f7, 'h100047, 'h100142, 'h10013e, 'h100143, 'h10013f, 'h100144, 'h100145, 'h100146, 'h100147, 'h100148, 'h100149, 'h10014a, 'h10014b, 'h10014c, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100140, 'h10003c, 'h2004f7, 'h100047, 'h100151, 'h10013d, 'h100152, 'h10013e, 'h100153, 'h10013f, 'h100154, 'h100155, 'h100156, 'h100157, 'h100158, 'h100159, 'h10015a, 'h10015b, 'h10015c, 'h10015e, 'h10015f, 'h100160, 'h10003c, 'h2004f7, 'h100047, 'h100140, 'h100162, 'h10013d, 'h10013e, 'h100163, 'h10013f, 'h100164, 'h100166, 'h100167, 'h100168, 'h10016a, 'h10016b, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h100145, 'h100144, 'h100147, 'h10003c, 'h2004f7, 'h100047, 'h100141, 'h100146, 'h100142, 'h100143, 'h100148, 'h100149, 'h10014b, 'h10014a, 'h10014c, 'h10014d, 'h10014f, 'h10014e, 'h100150, 'h100151, 'h100153, 'h100152, 'h100154, 'h100144, 'h10003c, 'h2004f7, 'h100047, 'h100155, 'h100157, 'h100156, 'h100141, 'h100142, 'h100143, 'h100158, 'h10015a, 'h10015b, 'h10015c, 'h10015e, 'h10015f, 'h100160, 'h100162, 'h100163, 'h100164, 'h100166, 'h100144, 'h100167, 'h10003c, 'h2004f7, 'h100047, 'h100168, 'h10016a, 'h10016b, 'h100141, 'h100142, 'h100143, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h100149, 'h100148, 'h10014a, 'h100145, 'h100146, 'h10014b, 'h100147, 'h10014c, 'h10003c, 'h2004f7, 'h100047, 'h10014d, 'h10014e, 'h10014f, 'h100150, 'h100151, 'h100152, 'h100153, 'h100154, 'h100156, 'h100157, 'h100158, 'h100148, 'h10015a, 'h100145, 'h100146, 'h10015b, 'h100147, 'h10015c, 'h10003c, 'h2004f7, 'h100047, 'h10015e, 'h10015f, 'h100160, 'h100162, 'h100163, 'h100164, 'h100166, 'h100167, 'h100168, 'h10016a, 'h10016b, 'h10016c, 'h100148, 'h10016e, 'h10016f, 'h100145, 'h100146, 'h100147, 'h10003c, 'h2004f7, 'h100047, 'h100170, 'h10014d, 'h10014c, 'h10014f, 'h10014e, 'h100149, 'h10014a, 'h10014b, 'h100150, 'h100152, 'h100153, 'h100154, 'h100156, 'h100157, 'h100158, 'h10015a, 'h10015b, 'h10015c, 'h10003c, 'h2004f7, 'h100047, 'h10015e, 'h10015f, 'h10014c, 'h100160, 'h100162, 'h100163, 'h100149, 'h10014a, 'h10014b, 'h100164, 'h100166, 'h100167, 'h100168, 'h10016a, 'h10016b, 'h10016c, 'h10016e, 'h10016f, 'h10003c, 'h2004f7, 'h100047, 'h100170, 'h100152, 'h100150, 'h10014e, 'h100153, 'h10014f, 'h100154, 'h100156, 'h100157, 'h100158, 'h10015a, 'h10015b, 'h10015c, 'h10015e, 'h10015f, 'h100160, 'h100162, 'h100163, 'h10003c, 'h2004f7, 'h100047, 'h100164, 'h100166, 'h100150, 'h10014e, 'h100167, 'h10014f, 'h100168, 'h10016a, 'h10016b, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h100156, 'h100154, 'h100152, 'h100157, 'h100153, 'h10003c, 'h2004f7, 'h100047, 'h100158, 'h10015a, 'h10015b, 'h10015c, 'h10015e, 'h10015f, 'h100160, 'h100162, 'h100163, 'h100164, 'h100166, 'h100167, 'h100168, 'h10016a, 'h100154, 'h100152, 'h10016b, 'h100153, 'h10003c, 'h2004f7, 'h100047, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h10015a, 'h100158, 'h100156, 'h10015b, 'h100157, 'h10015c, 'h10015e, 'h10015f, 'h100160, 'h100162, 'h100163, 'h100164, 'h100166, 'h100167, 'h10003c, 'h2004f7, 'h100047, 'h100168, 'h10016a, 'h10016b, 'h10016c, 'h10016e, 'h100158, 'h100156, 'h10016f, 'h100157, 'h100170, 'h10015e, 'h10015c, 'h10015a, 'h10015f, 'h10015b, 'h100160, 'h100162, 'h100163, 'h10003c, 'h2004f7, 'h100047, 'h100164, 'h100166, 'h100167, 'h100168, 'h10016a, 'h10016b, 'h10016c, 'h10016e, 'h10016f, 'h100170, 'h10015e, 'h2004f8, 'h100072, 'h100174, 'h10006e, 'h100171, 'h10006f, 'h100172, 'h100070, 'h10003c, 'h100047, 'h100173, 'h100071, 'h100178, 'h100175, 'h100176, 'h100177, 'h10017c, 'h100179, 'h10017a, 'h10017b, 'h100180, 'h2004f8, 'h100072, 'h10017d, 'h10006e, 'h10017e, 'h10006f, 'h10017f, 'h100070, 'h10003c, 'h100047, 'h100184, 'h100181, 'h100182, 'h100183, 'h100071, 'h100188, 'h100185, 'h100186, 'h100187, 'h10018c, 'h100189, 'h2004f8, 'h10018a, 'h10018b, 'h100072, 'h100190, 'h10006e, 'h10018d, 'h10006f, 'h10003c, 'h100047, 'h10018e, 'h100070, 'h10018f, 'h100194, 'h100191, 'h100192, 'h100193, 'h100071, 'h100198, 'h100195, 'h100196, 'h2004f8, 'h100197, 'h10019c, 'h100072, 'h100199, 'h10006e, 'h10019a, 'h10006f, 'h10003c, 'h100047, 'h10019b, 'h100070, 'h1001a0, 'h10019d, 'h10019e, 'h10019f, 'h1001a4, 'h1001a1, 'h1001a2, 'h1001a3, 'h100071, 'h2004f8, 'h1001a8, 'h1001a5, 'h1001a6, 'h1001a7, 'h100072, 'h1001a9, 'h1001ac, 'h10003c, 'h100047, 'h10006e, 'h10006f, 'h1001aa, 'h100070, 'h1001ab, 'h1001ad, 'h1001b0, 'h1001ae, 'h1001af, 'h1001b1, 'h1001b4, 'h2004f8, 'h1001b2, 'h1001b3, 'h100071, 'h1001b5, 'h100072, 'h1001b8, 'h1001b6, 'h10003c, 'h100047, 'h1001b7, 'h1001b9, 'h1001bc, 'h10006e, 'h10006f, 'h1001ba, 'h100070, 'h1001bb, 'h1001bd, 'h1001c0, 'h1001be, 'h2004f8, 'h1001bf, 'h1001c1, 'h1001c4, 'h1001c2, 'h1001c3, 'h100071, 'h100072, 'h10003c, 'h100047, 'h1001c5, 'h1001c8, 'h1001c6, 'h1001c7, 'h1001c9, 'h1001cc, 'h10006e, 'h10006f, 'h1001ca, 'h100070, 'h1001cb, 'h2004f8, 'h1001cd, 'h1001d0, 'h1001ce, 'h1001cf, 'h1001d1, 'h1001d4, 'h100072, 'h10003c, 'h100047, 'h1001d2, 'h1001d3, 'h100071, 'h1001d5, 'h1001d8, 'h1001d6, 'h1001d7, 'h1001d9, 'h1001dc, 'h10006e, 'h10006f, 'h2004f8, 'h1001da, 'h100070, 'h1001db, 'h1001dd, 'h1001e1, 'h1001de, 'h1001df, 'h10003c, 'h100047, 'h1001e0, 'h100072, 'h1001e5, 'h1001e2, 'h1001e3, 'h100071, 'h1001e4, 'h1001e9, 'h1001e6, 'h1001e7, 'h1001e8, 'h2004f8, 'h1001ed, 'h10006e, 'h10006f, 'h1001ea, 'h100070, 'h1001eb, 'h1001ec, 'h10003c, 'h100047, 'h1001f1, 'h100072, 'h1001ee, 'h1001ef, 'h1001f0, 'h100071, 'h1001f5, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f9, 'h2004f8, 'h1001f6, 'h10006e, 'h10006f, 'h1001f7, 'h100070, 'h1001f8, 'h1001fd, 'h10003c, 'h100047, 'h1001fa, 'h1001fb, 'h1001fc, 'h100072, 'h100201, 'h1001fe, 'h1001ff, 'h100200, 'h100071, 'h100205, 'h100202, 'h2004f8, 'h100203, 'h100204, 'h100209, 'h10006e, 'h100206, 'h10006f, 'h100207, 'h10003c, 'h100047, 'h100070, 'h100208, 'h10020d, 'h100072, 'h10020a, 'h10020b, 'h10020c, 'h100211, 'h10020e, 'h10020f, 'h100210, 'h2004f8, 'h100071, 'h100215, 'h100212, 'h10006e, 'h100213, 'h10006f, 'h100214, 'h10003c, 'h100047, 'h100070, 'h100219, 'h100216, 'h100217, 'h100218, 'h100072, 'h10021d, 'h10021a, 'h10021b, 'h10021c, 'h100221, 'h2004f8, 'h10021e, 'h10021f, 'h100220, 'h100071, 'h100225, 'h10006e, 'h100222, 'h10003c, 'h100047, 'h10006f, 'h100223, 'h100070, 'h100224, 'h100229, 'h100072, 'h100226, 'h100227, 'h100228, 'h10022a, 'h10022d, 'h2004f8, 'h10022b, 'h10022c, 'h10022e, 'h100231, 'h10022f, 'h100230, 'h100071, 'h10003c, 'h100047, 'h100232, 'h100235, 'h10006e, 'h10006f, 'h100233, 'h100070, 'h100234, 'h100072, 'h100236, 'h100239, 'h100237, 'h2004f8, 'h100238, 'h10023a, 'h10023d, 'h10023b, 'h10023c, 'h10023e, 'h100241, 'h10003c, 'h100047, 'h10023f, 'h100240, 'h100071, 'h100242, 'h100245, 'h10006e, 'h10006f, 'h100243, 'h100070, 'h100244, 'h100072, 'h2004f8, 'h100246, 'h100249, 'h100247, 'h100248, 'h10024a, 'h10024d, 'h10024b, 'h10003c, 'h100047, 'h10024c, 'h10024e, 'h100251, 'h10024f, 'h100250, 'h100071, 'h100252, 'h100255, 'h10006e, 'h10006f, 'h100253, 'h2004f8, 'h100070, 'h100254, 'h100072, 'h100256, 'h100259, 'h100257, 'h100258, 'h10003c, 'h100047, 'h10025a, 'h10025d, 'h10025b, 'h10025c, 'h10025e, 'h100262, 'h10025f, 'h100260, 'h100071, 'h100261, 'h100266, 'h2004f8, 'h10006e, 'h10006f, 'h100263, 'h100070, 'h100264, 'h100265, 'h100072, 'h10003c, 'h100047, 'h10026a, 'h100267, 'h100268, 'h100269, 'h10026e, 'h10026b, 'h10026c, 'h10026d, 'h100071, 'h100272, 'h10026f, 'h2004f8, 'h100270, 'h100271, 'h100170, 'h100076, 'h100073, 'h100171, 'h100074, 'h10003c, 'h100047, 'h100172, 'h100075, 'h100173, 'h100174, 'h100072, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h2004f8, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h100073, 'h10017f, 'h100074, 'h10003c, 'h100047, 'h100180, 'h100075, 'h100076, 'h100181, 'h100072, 'h100182, 'h100183, 'h100184, 'h100185, 'h100186, 'h100187, 'h2004f8, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h100073, 'h10003c, 'h100047, 'h10018e, 'h100074, 'h10018f, 'h100075, 'h100190, 'h100076, 'h100072, 'h100191, 'h100192, 'h100193, 'h100194, 'h2004f8, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h100073, 'h10003c, 'h100047, 'h10019b, 'h100074, 'h10019c, 'h100075, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h100076, 'h1001a1, 'h100072, 'h2004f8, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h10003c, 'h100047, 'h1001a9, 'h100073, 'h1001aa, 'h100074, 'h1001ab, 'h100075, 'h1001ac, 'h1001ad, 'h100076, 'h1001ae, 'h1001af, 'h2004f8, 'h1001b0, 'h1001b1, 'h100072, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h10003c, 'h100047, 'h1001b6, 'h100073, 'h1001b7, 'h100074, 'h1001b8, 'h100075, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h100076, 'h2004f8, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h100072, 'h1001c2, 'h10003c, 'h100047, 'h1001c3, 'h1001c4, 'h1001c5, 'h100073, 'h1001c6, 'h100074, 'h1001c7, 'h100075, 'h1001c8, 'h1001c9, 'h100076, 'h2004f8, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h10003c, 'h100047, 'h1001d1, 'h100072, 'h1001d2, 'h100073, 'h1001d3, 'h100074, 'h1001d4, 'h100075, 'h1001d5, 'h1001d6, 'h1001d7, 'h2004f8, 'h1001d8, 'h100076, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h10003c, 'h100047, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h100072, 'h100073, 'h1001e2, 'h100074, 'h1001e3, 'h100075, 'h1001e4, 'h2004f8, 'h1001e5, 'h100076, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h10003c, 'h100047, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h100072, 'h100073, 'h1001f2, 'h100074, 'h2004f8, 'h1001f3, 'h100075, 'h1001f4, 'h100076, 'h1001f5, 'h1001f6, 'h1001f7, 'h10003c, 'h100047, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h100072, 'h100073, 'h1001ff, 'h100074, 'h2004f8, 'h100200, 'h100075, 'h100201, 'h100076, 'h100202, 'h100203, 'h100204, 'h10003c, 'h100047, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h100072, 'h10020e, 'h2004f8, 'h100073, 'h10020f, 'h100074, 'h100210, 'h100075, 'h100211, 'h100076, 'h10003c, 'h100047, 'h100212, 'h100213, 'h100214, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h100072, 'h10021b, 'h2004f8, 'h100073, 'h10021c, 'h100074, 'h10021d, 'h100075, 'h10021e, 'h10021f, 'h10003c, 'h100047, 'h100220, 'h100221, 'h100076, 'h100222, 'h100223, 'h100224, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h2004f8, 'h10022a, 'h100072, 'h100073, 'h10022b, 'h100074, 'h10022c, 'h100075, 'h10003c, 'h100047, 'h10022d, 'h10022e, 'h100076, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h2004f8, 'h100237, 'h100238, 'h100239, 'h10023a, 'h100072, 'h100073, 'h10023b, 'h10003c, 'h100047, 'h100074, 'h10023c, 'h100075, 'h10023d, 'h100076, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h2004f8, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10003c, 'h100047, 'h100072, 'h100073, 'h10024b, 'h100074, 'h10024c, 'h100075, 'h10024d, 'h100076, 'h10024e, 'h10024f, 'h100250, 'h2004f8, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h10003c, 'h100047, 'h100258, 'h100259, 'h10025a, 'h100072, 'h100073, 'h10025b, 'h100074, 'h10025c, 'h100075, 'h10025d, 'h100076, 'h2004f8, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h10003c, 'h100047, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h100072, 'h100073, 'h10026b, 'h100074, 'h10026c, 'h2004f8, 'h100075, 'h10026d, 'h100076, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h10003c, 'h100047, 'h100272, 'h100170, 'h10007a, 'h100077, 'h100171, 'h100078, 'h100172, 'h100079, 'h100173, 'h100174, 'h100175, 'h2004f8, 'h100176, 'h100177, 'h100178, 'h100076, 'h100179, 'h10017a, 'h10017b, 'h10003c, 'h100047, 'h10017c, 'h10017d, 'h10017e, 'h100077, 'h10017f, 'h100078, 'h100180, 'h100079, 'h10007a, 'h100181, 'h100182, 'h2004f8, 'h100183, 'h100184, 'h100185, 'h100076, 'h100186, 'h100187, 'h100188, 'h10003c, 'h100047, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h100077, 'h10018e, 'h100078, 'h10018f, 'h100079, 'h100190, 'h2004f8, 'h10007a, 'h100191, 'h100192, 'h100193, 'h100194, 'h100076, 'h100195, 'h10003c, 'h100047, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h100077, 'h10019b, 'h100078, 'h10019c, 'h100079, 'h10019d, 'h2004f8, 'h10019e, 'h10019f, 'h1001a0, 'h10007a, 'h1001a1, 'h100076, 'h1001a2, 'h10003c, 'h100047, 'h1001a3, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h100077, 'h1001aa, 'h100078, 'h1001ab, 'h2004f8, 'h100079, 'h1001ac, 'h1001ad, 'h10007a, 'h1001ae, 'h1001af, 'h1001b0, 'h10003c, 'h100047, 'h1001b1, 'h100076, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h100077, 'h1001b7, 'h100078, 'h1001b8, 'h2004f8, 'h100079, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h10007a, 'h1001bd, 'h10003c, 'h100047, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h100076, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h100077, 'h1001c6, 'h2004f8, 'h100078, 'h1001c7, 'h100079, 'h1001c8, 'h1001c9, 'h10007a, 'h1001ca, 'h10003c, 'h100047, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h100076, 'h1001d2, 'h100077, 'h1001d3, 'h2004f8, 'h100078, 'h1001d4, 'h100079, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h10003c, 'h100047, 'h10007a, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h100076, 'h2004f8, 'h100077, 'h1001e2, 'h100078, 'h1001e3, 'h100079, 'h1001e4, 'h1001e5, 'h10003c, 'h100047, 'h10007a, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h2004f8, 'h1001f0, 'h1001f1, 'h100076, 'h100077, 'h1001f2, 'h100078, 'h1001f3, 'h10003c, 'h100047, 'h100079, 'h1001f4, 'h10007a, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h2004f8, 'h1001fd, 'h1001fe, 'h100076, 'h100077, 'h1001ff, 'h100078, 'h100200, 'h10003c, 'h100047, 'h100079, 'h100201, 'h10007a, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100207, 'h100208, 'h100209, 'h2004f8, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h100076, 'h10020e, 'h100077, 'h10003c, 'h100047, 'h10020f, 'h100078, 'h100210, 'h100079, 'h100211, 'h10007a, 'h100212, 'h100213, 'h100214, 'h100215, 'h100216, 'h2004f8, 'h100217, 'h100218, 'h100219, 'h10021a, 'h100076, 'h10021b, 'h100077, 'h10003c, 'h100047, 'h10021c, 'h100078, 'h10021d, 'h100079, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h10007a, 'h100222, 'h100223, 'h2004f8, 'h100224, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10003c, 'h100047, 'h100076, 'h100077, 'h10022b, 'h100078, 'h10022c, 'h100079, 'h10022d, 'h10022e, 'h10007a, 'h10022f, 'h100230, 'h2004f8, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h10003c, 'h100047, 'h100238, 'h100239, 'h10023a, 'h100076, 'h100077, 'h10023b, 'h100078, 'h10023c, 'h100079, 'h10023d, 'h10007a, 'h2004f8, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h10003c, 'h100047, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h100076, 'h100077, 'h10024b, 'h100078, 'h10024c, 'h2004f8, 'h100079, 'h10024d, 'h10007a, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h10003c, 'h100047, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h100076, 'h100077, 'h2004f8, 'h10025b, 'h100078, 'h10025c, 'h100079, 'h10025d, 'h10007a, 'h10025e, 'h10003c, 'h100047, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h2004f8, 'h10026a, 'h100076, 'h100077, 'h10026b, 'h100078, 'h10026c, 'h100079, 'h10003c, 'h100047, 'h10026d, 'h10007a, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100170, 'h10007e, 'h10007b, 'h100171, 'h2004f8, 'h10007c, 'h100172, 'h10007d, 'h100173, 'h100174, 'h100175, 'h100176, 'h10003c, 'h100047, 'h100177, 'h100178, 'h10007a, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h10007e, 'h2004f8, 'h100181, 'h10007b, 'h100182, 'h10007c, 'h100183, 'h10007d, 'h10003c, 'h100047, 'h100184, 'h100185, 'h10007a, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h2004f8, 'h10018f, 'h100190, 'h10007e, 'h100191, 'h10007b, 'h100192, 'h10003c, 'h100047, 'h10007c, 'h100193, 'h10007d, 'h100194, 'h10007a, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h2004f8, 'h10019c, 'h10019d, 'h10007e, 'h10019e, 'h10007b, 'h10019f, 'h10003c, 'h100047, 'h10007c, 'h1001a0, 'h10007d, 'h1001a1, 'h10007a, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h2004f8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h10007e, 'h1001ad, 'h10003c, 'h100047, 'h10007b, 'h1001ae, 'h10007c, 'h1001af, 'h10007d, 'h1001b0, 'h1001b1, 'h10007a, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h2004f8, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h10007e, 'h1001ba, 'h10003c, 'h100047, 'h10007b, 'h1001bb, 'h10007c, 'h1001bc, 'h10007d, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h10007a, 'h1001c2, 'h2004f8, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h10003c, 'h100047, 'h10007e, 'h1001c9, 'h10007b, 'h1001ca, 'h10007c, 'h1001cb, 'h10007d, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h2004f8, 'h1001d1, 'h10007a, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h10003c, 'h100047, 'h10007e, 'h1001d6, 'h10007b, 'h1001d7, 'h10007c, 'h1001d8, 'h10007d, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h2004f8, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h10007a, 'h1001e2, 'h10003c, 'h100047, 'h1001e3, 'h1001e4, 'h10007e, 'h1001e5, 'h10007b, 'h1001e6, 'h10007c, 'h1001e7, 'h10007d, 'h1001e8, 'h1001e9, 'h1001ea, 'h2004f8, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h10003c, 'h100047, 'h1001f1, 'h10007a, 'h1001f2, 'h1001f3, 'h1001f4, 'h10007e, 'h1001f5, 'h10007b, 'h1001f6, 'h10007c, 'h1001f7, 'h10007d, 'h2004f8, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h10003c, 'h100047, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h10007a, 'h100202, 'h100203, 'h10007b, 'h100204, 'h10007c, 'h100205, 'h10007d, 'h2004f8, 'h10007e, 'h100206, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10003c, 'h100047, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10007a, 'h10020f, 'h100210, 'h100211, 'h100212, 'h10007b, 'h100213, 'h10007c, 'h2004f8, 'h100214, 'h10007d, 'h100215, 'h10007e, 'h100216, 'h100217, 'h10003c, 'h100047, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10007a, 'h10021f, 'h10007b, 'h100220, 'h10007c, 'h2004f8, 'h100221, 'h10007d, 'h100222, 'h10007e, 'h100223, 'h100224, 'h10003c, 'h100047, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10007a, 'h10007b, 'h2004f8, 'h10022f, 'h10007c, 'h100230, 'h10007d, 'h100231, 'h10007e, 'h10003c, 'h100047, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h2004f8, 'h10023e, 'h10007a, 'h10007b, 'h10023f, 'h10007c, 'h100240, 'h10003c, 'h100047, 'h10007d, 'h100241, 'h10007e, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h2004f8, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10007a, 'h10007b, 'h10003c, 'h100047, 'h10024f, 'h10007c, 'h100250, 'h10007d, 'h100251, 'h10007e, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h2004f8, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10003c, 'h100047, 'h10025e, 'h10007a, 'h10007b, 'h10025f, 'h10007c, 'h100260, 'h10007d, 'h100261, 'h10007e, 'h100262, 'h100263, 'h100264, 'h2004f8, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10003c, 'h100047, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10007a, 'h10007b, 'h10026f, 'h10007c, 'h100270, 'h10007d, 'h100271, 'h10007e, 'h2004f8, 'h100272, 'h100170, 'h100082, 'h10007f, 'h100171, 'h100080, 'h10003c, 'h100047, 'h100172, 'h100081, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h2004f8, 'h10007e, 'h10017d, 'h10017e, 'h10017f, 'h100082, 'h100180, 'h10003c, 'h100047, 'h100181, 'h10007f, 'h100182, 'h100080, 'h100183, 'h100081, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h2004f8, 'h10007e, 'h10018a, 'h10018b, 'h10018c, 'h100082, 'h10018d, 'h10003c, 'h100047, 'h10018e, 'h10007f, 'h10018f, 'h100080, 'h100190, 'h100081, 'h100191, 'h100192, 'h100193, 'h100194, 'h100195, 'h100196, 'h2004f8, 'h100197, 'h100198, 'h100199, 'h10007e, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h10019c, 'h100082, 'h10019d, 'h10007f, 'h10019e, 'h100080, 'h10019f, 'h100081, 'h1001a0, 'h1001a1, 'h1001a2, 'h1001a3, 'h2004f8, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h10007e, 'h1001aa, 'h1001ab, 'h1001ac, 'h100082, 'h1001ad, 'h10007f, 'h1001ae, 'h100080, 'h1001af, 'h100081, 'h1001b0, 'h2004f8, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h10003c, 'h100047, 'h1001b7, 'h1001b8, 'h1001b9, 'h10007e, 'h1001ba, 'h1001bb, 'h1001bc, 'h100082, 'h1001bd, 'h10007f, 'h1001be, 'h100080, 'h2004f8, 'h1001bf, 'h100081, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h10003c, 'h100047, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h10007e, 'h1001ca, 'h1001cb, 'h1001cc, 'h100082, 'h1001cd, 'h2004f8, 'h10007f, 'h1001ce, 'h100080, 'h1001cf, 'h100081, 'h1001d0, 'h10003c, 'h100047, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h10007e, 'h1001da, 'h1001db, 'h2004f8, 'h1001dc, 'h100082, 'h1001dd, 'h10007f, 'h1001de, 'h100080, 'h10003c, 'h100047, 'h1001df, 'h100081, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h2004f8, 'h10007e, 'h1001ea, 'h1001eb, 'h1001ec, 'h100082, 'h1001ed, 'h10003c, 'h100047, 'h10007f, 'h1001ee, 'h100080, 'h1001ef, 'h100081, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h2004f8, 'h1001f7, 'h1001f8, 'h1001f9, 'h10007e, 'h1001fa, 'h1001fb, 'h10003c, 'h100047, 'h1001fc, 'h100082, 'h1001fd, 'h10007f, 'h1001fe, 'h100080, 'h1001ff, 'h100081, 'h100200, 'h100201, 'h100202, 'h100203, 'h2004f8, 'h100204, 'h100205, 'h100206, 'h10007e, 'h100207, 'h100208, 'h10003c, 'h100047, 'h100209, 'h100082, 'h10020a, 'h10007f, 'h10020b, 'h100080, 'h10020c, 'h100081, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h2004f8, 'h100211, 'h100212, 'h100213, 'h100214, 'h100215, 'h100216, 'h10007e, 'h10003c, 'h100047, 'h100217, 'h100218, 'h100219, 'h100082, 'h10021a, 'h10007f, 'h10021b, 'h100080, 'h10021c, 'h100081, 'h10021d, 'h2004f8, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h100223, 'h100224, 'h10003c, 'h100047, 'h100225, 'h100226, 'h10007e, 'h100227, 'h100228, 'h100229, 'h100082, 'h10022a, 'h10007f, 'h10022b, 'h100080, 'h2004f8, 'h10022c, 'h100081, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h10003c, 'h100047, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h10007e, 'h100237, 'h100238, 'h100239, 'h100082, 'h10023a, 'h2004f8, 'h10007f, 'h10023b, 'h100080, 'h10023c, 'h100081, 'h10023d, 'h10023e, 'h10003c, 'h100047, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h10007e, 'h100247, 'h100248, 'h2004f8, 'h100249, 'h100082, 'h10024a, 'h10007f, 'h10024b, 'h100080, 'h10024c, 'h10003c, 'h100047, 'h100081, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h2004f8, 'h10007e, 'h100257, 'h100258, 'h100259, 'h100082, 'h10025a, 'h10007f, 'h10003c, 'h100047, 'h10025b, 'h100080, 'h10025c, 'h100081, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h2004f8, 'h100264, 'h100265, 'h100266, 'h10007e, 'h100267, 'h100268, 'h100269, 'h10003c, 'h100047, 'h100082, 'h10026a, 'h10007f, 'h10026b, 'h100080, 'h10026c, 'h100081, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h2004f8, 'h100271, 'h100272, 'h100170, 'h100086, 'h100083, 'h100171, 'h100084, 'h10003c, 'h100047, 'h100172, 'h100085, 'h100173, 'h100174, 'h100082, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h2004f8, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100086, 'h100180, 'h10003c, 'h100047, 'h100083, 'h100181, 'h100084, 'h100182, 'h100085, 'h100183, 'h100184, 'h100082, 'h100185, 'h100186, 'h100187, 'h2004f8, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h100086, 'h10018d, 'h10003c, 'h100047, 'h100083, 'h10018e, 'h100084, 'h10018f, 'h100085, 'h100190, 'h100191, 'h100082, 'h100192, 'h100193, 'h100194, 'h2004f8, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h100086, 'h10019a, 'h10003c, 'h100047, 'h100083, 'h10019b, 'h100084, 'h10019c, 'h100085, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h100082, 'h2004f8, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h10003c, 'h100047, 'h100086, 'h1001a9, 'h100083, 'h1001aa, 'h100084, 'h1001ab, 'h100085, 'h1001ac, 'h1001ad, 'h1001ae, 'h1001af, 'h2004f8, 'h1001b0, 'h1001b1, 'h100082, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h10003c, 'h100047, 'h100086, 'h1001b6, 'h100083, 'h1001b7, 'h100084, 'h1001b8, 'h100085, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h2004f8, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h100082, 'h1001c2, 'h10003c, 'h100047, 'h1001c3, 'h1001c4, 'h100086, 'h1001c5, 'h100083, 'h1001c6, 'h100084, 'h1001c7, 'h100085, 'h1001c8, 'h1001c9, 'h2004f8, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h10003c, 'h100047, 'h1001d1, 'h100082, 'h1001d2, 'h1001d3, 'h1001d4, 'h100086, 'h1001d5, 'h100083, 'h1001d6, 'h100084, 'h1001d7, 'h2004f8, 'h100085, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h10003c, 'h100047, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h100082, 'h1001e2, 'h1001e3, 'h1001e4, 'h100086, 'h1001e5, 'h100083, 'h2004f8, 'h1001e6, 'h100084, 'h1001e7, 'h100085, 'h1001e8, 'h1001e9, 'h1001ea, 'h10003c, 'h100047, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h100082, 'h1001f2, 'h1001f3, 'h1001f4, 'h2004f8, 'h100086, 'h1001f5, 'h100083, 'h1001f6, 'h100084, 'h1001f7, 'h100085, 'h10003c, 'h100047, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100082, 'h2004f8, 'h100202, 'h100203, 'h100204, 'h100086, 'h100205, 'h100206, 'h100083, 'h10003c, 'h100047, 'h100207, 'h100084, 'h100208, 'h100085, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h100082, 'h2004f8, 'h10020f, 'h100210, 'h100211, 'h100086, 'h100212, 'h100213, 'h100083, 'h10003c, 'h100047, 'h100214, 'h100084, 'h100215, 'h100085, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h2004f8, 'h10021d, 'h10021e, 'h100082, 'h10021f, 'h100220, 'h100221, 'h100086, 'h10003c, 'h100047, 'h100222, 'h100083, 'h100223, 'h100084, 'h100224, 'h100085, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h2004f8, 'h10022a, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h100082, 'h10022f, 'h10003c, 'h100047, 'h100230, 'h100231, 'h100086, 'h100232, 'h100083, 'h100233, 'h100084, 'h100234, 'h100085, 'h100235, 'h100236, 'h2004f8, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10003c, 'h100047, 'h10023e, 'h100082, 'h10023f, 'h100240, 'h100241, 'h100086, 'h100242, 'h100083, 'h100243, 'h100084, 'h100244, 'h2004f8, 'h100085, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10003c, 'h100047, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h100082, 'h10024f, 'h100250, 'h100251, 'h100086, 'h100252, 'h100083, 'h2004f8, 'h100253, 'h100084, 'h100254, 'h100085, 'h100255, 'h100256, 'h100257, 'h10003c, 'h100047, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h100082, 'h10025f, 'h100260, 'h100261, 'h2004f8, 'h100086, 'h100262, 'h100083, 'h100263, 'h100084, 'h100264, 'h100085, 'h10003c, 'h100047, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h100082, 'h2004f8, 'h10026f, 'h100270, 'h100271, 'h100086, 'h100272, 'h100170, 'h10008a, 'h10003c, 'h100047, 'h100087, 'h100171, 'h100088, 'h100172, 'h100089, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h2004f8, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h100086, 'h10017d, 'h10017e, 'h10003c, 'h100047, 'h10017f, 'h10008a, 'h100180, 'h100087, 'h100181, 'h100088, 'h100182, 'h100089, 'h100183, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10003c, 'h100047, 'h10018d, 'h100086, 'h10018e, 'h100087, 'h10018f, 'h100088, 'h100190, 'h100089, 'h10008a, 'h100191, 'h100192, 'h2004f8, 'h100193, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10003c, 'h100047, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h100086, 'h100087, 'h10019e, 'h100088, 'h10019f, 'h100089, 'h1001a0, 'h2004f8, 'h10008a, 'h1001a1, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a5, 'h1001a6, 'h10003c, 'h100047, 'h1001a7, 'h1001a8, 'h1001a9, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ad, 'h100086, 'h100087, 'h1001ae, 'h100088, 'h2004f8, 'h1001af, 'h100089, 'h1001b0, 'h10008a, 'h1001b1, 'h1001b2, 'h1001b3, 'h10003c, 'h100047, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h100086, 'h2004f8, 'h100087, 'h1001be, 'h100088, 'h1001bf, 'h100089, 'h1001c0, 'h10008a, 'h10003c, 'h100047, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h2004f8, 'h1001cc, 'h1001cd, 'h100086, 'h100087, 'h1001ce, 'h100088, 'h1001cf, 'h10003c, 'h100047, 'h100089, 'h1001d0, 'h10008a, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h2004f8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h100086, 'h100087, 'h10003c, 'h100047, 'h1001de, 'h100088, 'h1001df, 'h100089, 'h1001e0, 'h10008a, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h2004f8, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h10003c, 'h100047, 'h1001ed, 'h100086, 'h100087, 'h1001ee, 'h100088, 'h1001ef, 'h100089, 'h1001f0, 'h10008a, 'h1001f1, 'h1001f2, 'h2004f8, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h10003c, 'h100047, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h100086, 'h100087, 'h1001fe, 'h100088, 'h1001ff, 'h100089, 'h100200, 'h2004f8, 'h10008a, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h10003c, 'h100047, 'h100207, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h100086, 'h100087, 'h10020f, 'h2004f8, 'h100088, 'h100210, 'h100089, 'h100211, 'h10008a, 'h100212, 'h100213, 'h10003c, 'h100047, 'h100214, 'h100215, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h2004f8, 'h100086, 'h100087, 'h10021f, 'h100088, 'h100220, 'h100089, 'h100221, 'h10003c, 'h100047, 'h10008a, 'h100222, 'h100223, 'h100224, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10022b, 'h2004f8, 'h10022c, 'h10022d, 'h10022e, 'h100086, 'h100087, 'h10022f, 'h100088, 'h10003c, 'h100047, 'h100230, 'h100089, 'h100231, 'h10008a, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h2004f8, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h100086, 'h10003c, 'h100047, 'h100087, 'h10023f, 'h100088, 'h100240, 'h100089, 'h100241, 'h10008a, 'h100242, 'h100243, 'h100244, 'h100245, 'h2004f8, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10003c, 'h100047, 'h10024d, 'h10024e, 'h100086, 'h100087, 'h10024f, 'h100088, 'h100250, 'h100089, 'h100251, 'h10008a, 'h100252, 'h2004f8, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10003c, 'h100047, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h100086, 'h100087, 'h10025f, 'h100088, 'h100260, 'h100089, 'h2004f8, 'h100261, 'h10008a, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h10003c, 'h100047, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h100086, 'h100087, 'h10026f, 'h2004f8, 'h100088, 'h100270, 'h100089, 'h100271, 'h10008a, 'h100272, 'h100170, 'h10008e, 'h10003c, 'h100047, 'h10008b, 'h100171, 'h10008c, 'h100172, 'h10008d, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h2004f8, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h10008e, 'h100180, 'h10008b, 'h100181, 'h10008c, 'h100182, 'h10008d, 'h100183, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h10008e, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h10008b, 'h100192, 'h10008c, 'h100193, 'h10008d, 'h2004f8, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h10019c, 'h10008e, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h10008b, 'h1001a2, 'h10008c, 'h2004f8, 'h1001a3, 'h10008d, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h1001aa, 'h1001ab, 'h1001ac, 'h10008e, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h10008b, 'h2004f8, 'h1001b2, 'h10008c, 'h1001b3, 'h10008d, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h100047, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h10008e, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h2004f8, 'h1001c1, 'h10008b, 'h1001c2, 'h10008c, 'h1001c3, 'h10008d, 'h1001c4, 'h1001c5, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h10008e, 'h1001cd, 'h1001ce, 'h2004f8, 'h1001cf, 'h1001d0, 'h1001d1, 'h10008b, 'h1001d2, 'h10008c, 'h1001d3, 'h10008d, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h10008e, 'h2004f8, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h10008b, 'h1001e2, 'h10008c, 'h10003c, 'h100047, 'h1001e3, 'h10008d, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h2004f8, 'h1001ec, 'h10008e, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h10008b, 'h10003c, 'h100047, 'h1001f2, 'h10008c, 'h1001f3, 'h10008d, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h2004f8, 'h1001fa, 'h1001fb, 'h1001fc, 'h10008e, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h10003c, 'h100047, 'h100201, 'h10008b, 'h100202, 'h10008c, 'h100203, 'h10008d, 'h100204, 'h100205, 'h100206, 'h100207, 'h2004f8, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10008e, 'h10020d, 'h10020e, 'h10003c, 'h100047, 'h10020f, 'h100210, 'h100211, 'h100212, 'h10008b, 'h100213, 'h10008c, 'h100214, 'h10008d, 'h100215, 'h2004f8, 'h100216, 'h100217, 'h100218, 'h100219, 'h10021a, 'h10008e, 'h10021b, 'h10021c, 'h10003c, 'h100047, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h10008b, 'h100223, 'h10008c, 'h100224, 'h2004f8, 'h10008d, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h10008e, 'h10022a, 'h10003c, 'h100047, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h10008b, 'h100233, 'h2004f8, 'h10008c, 'h100234, 'h10008d, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10003c, 'h100047, 'h10008e, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h2004f8, 'h10008b, 'h100243, 'h10008c, 'h100244, 'h10008d, 'h100245, 'h100246, 'h100247, 'h10003c, 'h100047, 'h100248, 'h100249, 'h10008e, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h2004f8, 'h100251, 'h100252, 'h10008b, 'h100253, 'h10008c, 'h100254, 'h10008d, 'h100255, 'h10003c, 'h100047, 'h100256, 'h100257, 'h100258, 'h100259, 'h10008e, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h2004f8, 'h10025f, 'h100260, 'h100261, 'h100262, 'h10008b, 'h100263, 'h10008c, 'h100264, 'h10003c, 'h100047, 'h10008d, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10008e, 'h10026a, 'h10026b, 'h10026c, 'h2004f8, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100170, 'h100092, 'h10003c, 'h100047, 'h10008f, 'h100171, 'h100090, 'h100172, 'h100091, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h2004f8, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h100092, 'h100180, 'h10008f, 'h100181, 'h100090, 'h100182, 'h100091, 'h100183, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h100092, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h10008f, 'h100192, 'h100090, 'h100193, 'h100091, 'h2004f8, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h10019c, 'h100092, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h10008f, 'h1001a2, 'h100090, 'h2004f8, 'h1001a3, 'h100091, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h1001aa, 'h1001ab, 'h1001ac, 'h100092, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h10008f, 'h2004f8, 'h1001b2, 'h100090, 'h1001b3, 'h100091, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h100047, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h100092, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h2004f8, 'h1001c1, 'h10008f, 'h1001c2, 'h100090, 'h1001c3, 'h100091, 'h1001c4, 'h1001c5, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h100092, 'h1001cd, 'h1001ce, 'h2004f8, 'h1001cf, 'h1001d0, 'h1001d1, 'h10008f, 'h1001d2, 'h100090, 'h1001d3, 'h100091, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h100092, 'h2004f8, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h10008f, 'h1001e2, 'h100090, 'h10003c, 'h100047, 'h1001e3, 'h100091, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h2004f8, 'h1001ec, 'h100092, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h10008f, 'h10003c, 'h100047, 'h1001f2, 'h100090, 'h1001f3, 'h100091, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h2004f8, 'h1001fa, 'h1001fb, 'h1001fc, 'h100092, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h10003c, 'h100047, 'h100201, 'h10008f, 'h100202, 'h100090, 'h100203, 'h100091, 'h100204, 'h100205, 'h100206, 'h100207, 'h2004f8, 'h100208, 'h100209, 'h10020a, 'h100092, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10003c, 'h100047, 'h10020f, 'h100210, 'h100211, 'h100212, 'h10008f, 'h100213, 'h100090, 'h100214, 'h100091, 'h100215, 'h2004f8, 'h100216, 'h100217, 'h100218, 'h100219, 'h100092, 'h10021a, 'h10021b, 'h10021c, 'h10003c, 'h100047, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h10008f, 'h100223, 'h100090, 'h100224, 'h2004f8, 'h100091, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h100092, 'h10022a, 'h10003c, 'h100047, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h10008f, 'h100233, 'h2004f8, 'h100090, 'h100234, 'h100091, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10003c, 'h100047, 'h100092, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h2004f8, 'h10008f, 'h100243, 'h100090, 'h100244, 'h100091, 'h100245, 'h100246, 'h100247, 'h10003c, 'h100047, 'h100248, 'h100249, 'h100092, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h2004f8, 'h100251, 'h100252, 'h10008f, 'h100253, 'h100090, 'h100254, 'h100091, 'h100255, 'h10003c, 'h100047, 'h100256, 'h100257, 'h100258, 'h100259, 'h100092, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h2004f8, 'h10025f, 'h100260, 'h100261, 'h100262, 'h10008f, 'h100263, 'h100090, 'h100264, 'h10003c, 'h100047, 'h100091, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h100092, 'h10026a, 'h10026b, 'h10026c, 'h2004f8, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100170, 'h100096, 'h10003c, 'h100047, 'h100093, 'h100171, 'h100094, 'h100172, 'h100095, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h2004f8, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h100096, 'h100180, 'h100181, 'h100093, 'h100094, 'h100182, 'h100095, 'h100183, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h100096, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h100093, 'h100094, 'h100192, 'h100095, 'h100193, 'h2004f8, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h10019c, 'h100096, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h100093, 'h1001a2, 'h100094, 'h2004f8, 'h1001a3, 'h100095, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h1001aa, 'h1001ab, 'h1001ac, 'h100096, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h100093, 'h2004f8, 'h1001b2, 'h100094, 'h1001b3, 'h100095, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h100047, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h100096, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h2004f8, 'h1001c1, 'h100093, 'h1001c2, 'h100094, 'h1001c3, 'h100095, 'h1001c4, 'h1001c5, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h100096, 'h1001cd, 'h1001ce, 'h2004f8, 'h1001cf, 'h1001d0, 'h1001d1, 'h100093, 'h1001d2, 'h100094, 'h1001d3, 'h100095, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h100096, 'h2004f8, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h100093, 'h1001e2, 'h100094, 'h10003c, 'h100047, 'h1001e3, 'h100095, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h2004f8, 'h1001ec, 'h100096, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h100093, 'h10003c, 'h100047, 'h1001f2, 'h100094, 'h1001f3, 'h100095, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h2004f8, 'h1001fa, 'h1001fb, 'h1001fc, 'h100096, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h10003c, 'h100047, 'h100201, 'h100202, 'h100093, 'h100094, 'h100203, 'h100095, 'h100204, 'h100205, 'h100206, 'h100207, 'h2004f8, 'h100208, 'h100209, 'h10020a, 'h100096, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10003c, 'h100047, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100093, 'h100094, 'h100213, 'h100095, 'h100214, 'h100215, 'h2004f8, 'h100216, 'h100217, 'h100218, 'h100219, 'h100096, 'h10021a, 'h10021b, 'h10021c, 'h10003c, 'h100047, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h100093, 'h100223, 'h100094, 'h100224, 'h2004f8, 'h100095, 'h100225, 'h100226, 'h100227, 'h100228, 'h100229, 'h100096, 'h10022a, 'h10003c, 'h100047, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100093, 'h100233, 'h2004f8, 'h100094, 'h100234, 'h100095, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10003c, 'h100047, 'h100096, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h2004f8, 'h100093, 'h100243, 'h100094, 'h100244, 'h100095, 'h100245, 'h100246, 'h100247, 'h10003c, 'h100047, 'h100248, 'h100249, 'h100096, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h2004f8, 'h100251, 'h100252, 'h100093, 'h100253, 'h100094, 'h100254, 'h100095, 'h100255, 'h10003c, 'h100047, 'h100256, 'h100257, 'h100258, 'h100259, 'h100096, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h2004f8, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100093, 'h100263, 'h100094, 'h100264, 'h10003c, 'h100047, 'h100095, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h100096, 'h10026a, 'h10026b, 'h10026c, 'h2004f8, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100170, 'h10009a, 'h10003c, 'h100047, 'h100097, 'h100171, 'h100098, 'h100172, 'h100099, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h2004f8, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10003c, 'h100047, 'h10009a, 'h100180, 'h100181, 'h100097, 'h100098, 'h100182, 'h100099, 'h100183, 'h100184, 'h100185, 'h2004f8, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10003c, 'h100047, 'h10009a, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h100097, 'h100098, 'h100192, 'h100099, 'h100193, 'h2004f8, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10003c, 'h100047, 'h10019c, 'h10009a, 'h10019d, 'h10019e, 'h10019f, 'h1001a0, 'h1001a1, 'h100097, 'h1001a2, 'h100098, 'h2004f8, 'h1001a3, 'h100099, 'h1001a4, 'h1001a5, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001a9, 'h10003c, 'h100047, 'h1001aa, 'h1001ab, 'h1001ac, 'h10009a, 'h1001ad, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h100097, 'h2004f8, 'h1001b2, 'h100098, 'h1001b3, 'h100099, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h100047, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h10009a, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h2004f8, 'h1001c1, 'h100097, 'h1001c2, 'h100098, 'h1001c3, 'h100099, 'h1001c4, 'h1001c5, 'h10003c, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h10009a, 'h1001cd, 'h1001ce, 'h2004f8, 'h1001cf, 'h1001d0, 'h1001d1, 'h100097, 'h1001d2, 'h100098, 'h1001d3, 'h100099, 'h10003c, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h10009a, 'h2004f8, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h100097, 'h1001e2, 'h100098, 'h10003c, 'h100047, 'h1001e3, 'h100099, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h2004f8, 'h1001ec, 'h10009a, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h100097, 'h10003c, 'h100047, 'h1001f2, 'h100098, 'h1001f3, 'h100099, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h1001f9, 'h2004f8, 'h1001fa, 'h1001fb, 'h1001fc, 'h10009a, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h10003c, 'h100047, 'h100201, 'h100202, 'h100097, 'h100098, 'h100203, 'h100099, 'h100204, 'h100205, 'h100206, 'h100207, 'h2004f8, 'h100208, 'h100209, 'h10020a, 'h10009a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10003c, 'h100047, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100097, 'h100098, 'h100213, 'h100099, 'h100214, 'h100215, 'h2004f8, 'h100216, 'h100217, 'h100218, 'h10009a, 'h100219, 'h10021a, 'h10021b, 'h10021c, 'h10003c, 'h100047, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h100222, 'h100097, 'h100223, 'h100098, 'h100224, 'h2004f8, 'h100099, 'h100225, 'h100226, 'h10009a, 'h100227, 'h100228, 'h100229, 'h10022a, 'h10003c, 'h100047, 'h10022b, 'h10022c, 'h10022d, 'h10022e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100097, 'h100233, 'h2004f8, 'h100098, 'h100234, 'h100099, 'h100235, 'h10009a, 'h100236, 'h100237, 'h100238, 'h10003c, 'h100047, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h2004f8, 'h100097, 'h100243, 'h100098, 'h100244, 'h100099, 'h100245, 'h10009a, 'h100246, 'h10003c, 'h100047, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h2004f8, 'h100251, 'h100252, 'h100097, 'h100253, 'h100098, 'h100254, 'h100099, 'h100255, 'h10003c, 'h100047, 'h10009a, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h2004f8, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100097, 'h100263, 'h100098, 'h100264, 'h10003c, 'h100047, 'h100099, 'h100265, 'h10009a, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b};
	int DATA2 [2*SIZE-1:0] = {DATA1, DATA0};
	
endpackage
