

package MATRIX_MULTIPLY_32_PKG_1;
	
	parameter SIZE = 8500;
	
	int DATA1 [SIZE-1:0] = {'h21f91, 'h103be, 'h106b8, 'h21f90, 'h21f8f, 'h21f8d, 'h103c0, 'h21f8a, 'h21f8c, 'h103c1, 'h11f9c, 'h103bc, 'h10005, 'h11f9d, 'h10002, 'h21f8e, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106de, 'h106df, 'h106e0, 'h21f8c, 'h106e1, 'h106e2, 'h103bc, 'h106e3, 'h106e4, 'h106e5, 'h106e6, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h106e7, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106e8, 'h106e9, 'h21f8c, 'h106ea, 'h106eb, 'h103bc, 'h106ec, 'h106ed, 'h106ee, 'h106ef, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h106f0, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106f1, 'h106f2, 'h21f8c, 'h106f3, 'h106f4, 'h103bc, 'h106f5, 'h106f6, 'h106f7, 'h106f8, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h106f9, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106fa, 'h106fb, 'h21f8c, 'h106fc, 'h106fd, 'h103bc, 'h106fe, 'h106ff, 'h10700, 'h10701, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10702, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10703, 'h10704, 'h21f8c, 'h10705, 'h10706, 'h103bc, 'h10707, 'h10708, 'h10709, 'h1070a, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1070b, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1070c, 'h1070d, 'h21f8c, 'h1070e, 'h1070f, 'h103bc, 'h10710, 'h10711, 'h10712, 'h10713, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10714, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10715, 'h10716, 'h21f8c, 'h10717, 'h10718, 'h103bc, 'h10719, 'h1071a, 'h1071b, 'h1071c, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1071d, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1071e, 'h1071f, 'h21f8c, 'h10720, 'h10721, 'h103bc, 'h10722, 'h10723, 'h10724, 'h10725, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10726, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10727, 'h10728, 'h21f8c, 'h10729, 'h1072a, 'h103bc, 'h1072b, 'h1072c, 'h1072d, 'h1072e, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1072f, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10730, 'h10731, 'h21f8c, 'h10732, 'h10733, 'h103bc, 'h10734, 'h10735, 'h10736, 'h10737, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10738, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10739, 'h1073a, 'h21f8c, 'h1073b, 'h1073c, 'h103bc, 'h1073d, 'h1073e, 'h1073f, 'h10740, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10741, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10742, 'h10743, 'h21f8c, 'h10744, 'h10745, 'h103bc, 'h10746, 'h10747, 'h10748, 'h10749, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1074a, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1074b, 'h1074c, 'h21f8c, 'h1074d, 'h1074e, 'h103bc, 'h1074f, 'h10750, 'h10751, 'h10752, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10753, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10754, 'h10755, 'h21f8c, 'h10756, 'h10757, 'h103bc, 'h10758, 'h10759, 'h1075a, 'h1075b, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1075c, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1075d, 'h1075e, 'h21f8c, 'h1075f, 'h10760, 'h103bc, 'h10761, 'h10762, 'h10763, 'h10764, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10765, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10766, 'h10767, 'h21f8c, 'h10768, 'h10769, 'h103bc, 'h1076a, 'h1076b, 'h1076c, 'h1076d, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1076e, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1076f, 'h10770, 'h21f8c, 'h10771, 'h10772, 'h103bc, 'h10773, 'h10774, 'h10775, 'h10776, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10777, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10778, 'h10779, 'h21f8c, 'h1077a, 'h1077b, 'h103bc, 'h1077c, 'h1077d, 'h1077e, 'h1077f, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10780, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10781, 'h10782, 'h21f8c, 'h10783, 'h10784, 'h103bc, 'h10785, 'h10786, 'h10787, 'h10788, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10789, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1078a, 'h1078b, 'h21f8c, 'h1078c, 'h1078d, 'h103bc, 'h1078e, 'h1078f, 'h10790, 'h10791, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10792, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10793, 'h10794, 'h21f8c, 'h10795, 'h10796, 'h103bc, 'h10797, 'h10798, 'h10799, 'h1079a, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1079b, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1079c, 'h1079d, 'h21f8c, 'h1079e, 'h1079f, 'h103bc, 'h107a0, 'h107a1, 'h107a2, 'h107a3, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107a4, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107a5, 'h107a6, 'h21f8c, 'h107a7, 'h107a8, 'h103bc, 'h107a9, 'h107aa, 'h107ab, 'h107ac, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107ad, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107ae, 'h107af, 'h21f8c, 'h107b0, 'h107b1, 'h103bc, 'h107b2, 'h107b3, 'h107b4, 'h107b5, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107b6, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107b7, 'h107b8, 'h21f8c, 'h107b9, 'h107ba, 'h103bc, 'h107bb, 'h107bc, 'h107bd, 'h107be, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107c0, 'h107c1, 'h21f8c, 'h107c2, 'h107c3, 'h103bc, 'h107c4, 'h107c5, 'h107c6, 'h107c7, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107c8, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107c9, 'h107ca, 'h21f8c, 'h107cb, 'h107cc, 'h103bc, 'h107cd, 'h107ce, 'h107cf, 'h107d0, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107d1, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107d2, 'h107d3, 'h21f8c, 'h107d4, 'h107d5, 'h103bc, 'h107d6, 'h107d7, 'h107d8, 'h107d9, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107da, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107db, 'h107dc, 'h21f8c, 'h107dd, 'h107de, 'h103bc, 'h107df, 'h107e0, 'h107e1, 'h107e2, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107e3, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107e4, 'h107e5, 'h21f8c, 'h107e6, 'h107e7, 'h103bc, 'h107e8, 'h107e9, 'h107ea, 'h107eb, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107ec, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107ed, 'h107ee, 'h21f8c, 'h107ef, 'h107f0, 'h103bc, 'h107f1, 'h107f2, 'h107f3, 'h107f4, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107f5, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107f6, 'h107f7, 'h21f8c, 'h107f8, 'h107f9, 'h103bc, 'h107fa, 'h107fb, 'h107fc, 'h107fd, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107fe, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107ff, 'h10800, 'h21f8c, 'h10801, 'h10802, 'h103bc, 'h10803, 'h10804, 'h10805, 'h10806, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10807, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10808, 'h10809, 'h21f8c, 'h1080a, 'h1080b, 'h103bc, 'h1080c, 'h1080d, 'h1080e, 'h1080f, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10810, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10811, 'h10812, 'h21f8c, 'h10813, 'h10814, 'h103bc, 'h10815, 'h10816, 'h10817, 'h10818, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10819, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1081a, 'h1081b, 'h21f8c, 'h1081c, 'h1081d, 'h103bc, 'h1081e, 'h1081f, 'h10820, 'h10821, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10822, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10823, 'h10824, 'h21f8c, 'h10825, 'h10826, 'h103bc, 'h10827, 'h10828, 'h10829, 'h1082a, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1082b, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1082c, 'h1082d, 'h21f8c, 'h1082e, 'h1082f, 'h103bc, 'h10830, 'h10831, 'h10832, 'h10833, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10834, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10835, 'h10836, 'h21f8c, 'h10837, 'h10838, 'h103bc, 'h10839, 'h1083a, 'h1083b, 'h1083c, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1083d, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1083e, 'h1083f, 'h21f8c, 'h10840, 'h10841, 'h103bc, 'h10842, 'h10843, 'h10844, 'h10845, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10846, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10847, 'h10848, 'h21f8c, 'h10849, 'h1084a, 'h103bc, 'h1084b, 'h1084c, 'h1084d, 'h1084e, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1084f, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10850, 'h10851, 'h21f8c, 'h10852, 'h10853, 'h103bc, 'h10854, 'h10855, 'h10856, 'h10857, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10858, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10859, 'h1085a, 'h21f8c, 'h1085b, 'h1085c, 'h103bc, 'h1085d, 'h1085e, 'h1085f, 'h10860, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10861, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10862, 'h10863, 'h21f8c, 'h10864, 'h10865, 'h103bc, 'h10866, 'h10867, 'h10868, 'h10869, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1086a, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1086b, 'h1086c, 'h21f8c, 'h1086d, 'h1086e, 'h103bc, 'h1086f, 'h10870, 'h10871, 'h10872, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10873, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10874, 'h10875, 'h21f8c, 'h10876, 'h10877, 'h103bc, 'h10878, 'h10879, 'h1087a, 'h1087b, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1087c, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1087d, 'h1087e, 'h21f8c, 'h1087f, 'h10880, 'h103bc, 'h10881, 'h10882, 'h10883, 'h10884, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10885, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10886, 'h10887, 'h21f8c, 'h10888, 'h10889, 'h103bc, 'h1088a, 'h1088b, 'h1088c, 'h1088d, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1088e, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1088f, 'h10890, 'h21f8c, 'h10891, 'h10892, 'h103bc, 'h10893, 'h10894, 'h10895, 'h10896, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10897, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10898, 'h10899, 'h21f8c, 'h1089a, 'h1089b, 'h103bc, 'h1089c, 'h1089d, 'h1089e, 'h1089f, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h108a0, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108a1, 'h108a2, 'h21f8c, 'h108a3, 'h108a4, 'h103bc, 'h108a5, 'h108a6, 'h108a7, 'h108a8, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h108a9, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108aa, 'h108ab, 'h21f8c, 'h108ac, 'h108ad, 'h103bc, 'h108ae, 'h108af, 'h108b0, 'h108b1, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h108b2, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108b3, 'h108b4, 'h21f8c, 'h108b5, 'h108b6, 'h103bc, 'h108b7, 'h108b8, 'h108b9, 'h108ba, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h108bb, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108bc, 'h108bd, 'h21f8c, 'h108be, 'h108bf, 'h103bc, 'h108c0, 'h108c1, 'h108c2, 'h108c3, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h108c4, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108c5, 'h108c6, 'h21f8c, 'h108c7, 'h108c8, 'h103bc, 'h108c9, 'h108ca, 'h108cb, 'h108cc, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h108cd, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108ce, 'h108cf, 'h21f8c, 'h108d0, 'h108d1, 'h103bc, 'h108d2, 'h108d3, 'h108d4, 'h108d5, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h108d6, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108d7, 'h108d8, 'h21f8c, 'h108d9, 'h108da, 'h103bc, 'h108db, 'h108dc, 'h108dd, 'h21f8d, 'h10001, 'h10000, 'h108de, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108df, 'h108e0, 'h21f8c, 'h108e1, 'h108e2, 'h103bc, 'h108e3, 'h108e4, 'h108e5, 'h108e6, 'h10001, 'h10000, 'h108e7, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108e8, 'h108e9, 'h21f8c, 'h108ea, 'h108eb, 'h103bc, 'h108ec, 'h108ed, 'h108ee, 'h108ef, 'h10001, 'h10000, 'h108f0, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108f1, 'h108f2, 'h21f8c, 'h108f3, 'h108f4, 'h103bc, 'h108f5, 'h108f6, 'h108f7, 'h108f8, 'h10001, 'h10000, 'h108f9, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h108fa, 'h108fb, 'h21f8c, 'h108fc, 'h108fd, 'h103bc, 'h108fe, 'h108ff, 'h10900, 'h10901, 'h10001, 'h10000, 'h10902, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10903, 'h10904, 'h21f8c, 'h10905, 'h10906, 'h103bc, 'h10907, 'h10908, 'h10909, 'h1090a, 'h10001, 'h10000, 'h1090b, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1090c, 'h1090d, 'h21f8c, 'h1090e, 'h1090f, 'h103bc, 'h10910, 'h10911, 'h10912, 'h10913, 'h10001, 'h10000, 'h10914, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10915, 'h10916, 'h21f8c, 'h10917, 'h10918, 'h103bc, 'h10919, 'h1091a, 'h1091b, 'h1091c, 'h10001, 'h10000, 'h1091d, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1091e, 'h1091f, 'h21f8c, 'h10920, 'h10921, 'h103bc, 'h10922, 'h10923, 'h10924, 'h10925, 'h10001, 'h10000, 'h10926, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10927, 'h10928, 'h21f8c, 'h10929, 'h1092a, 'h103bc, 'h1092b, 'h1092c, 'h1092d, 'h1092e, 'h10001, 'h10000, 'h1092f, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10930, 'h10931, 'h21f8c, 'h10932, 'h10933, 'h103bc, 'h10934, 'h10935, 'h10936, 'h10937, 'h10001, 'h10000, 'h10938, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10939, 'h1093a, 'h21f8c, 'h1093b, 'h1093c, 'h103bc, 'h1093d, 'h1093e, 'h1093f, 'h10940, 'h10001, 'h10000, 'h10941, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10942, 'h10943, 'h21f8c, 'h10944, 'h10945, 'h103bc, 'h10946, 'h10947, 'h10948, 'h10949, 'h10001, 'h10000, 'h1094a, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1094b, 'h1094c, 'h21f8c, 'h1094d, 'h1094e, 'h103bc, 'h1094f, 'h10950, 'h10951, 'h10952, 'h10001, 'h10000, 'h10953, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10954, 'h10955, 'h21f8c, 'h10956, 'h10957, 'h103bc, 'h10958, 'h10959, 'h1095a, 'h1095b, 'h10001, 'h10000, 'h1095c, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1095d, 'h1095e, 'h21f8c, 'h1095f, 'h10960, 'h103bc, 'h10961, 'h10962, 'h10963, 'h10964, 'h10001, 'h10000, 'h10965, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10966, 'h10967, 'h21f8c, 'h10968, 'h10969, 'h103bc, 'h1096a, 'h1096b, 'h1096c, 'h1096d, 'h10001, 'h10000, 'h1096e, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1096f, 'h10970, 'h21f8c, 'h10971, 'h10972, 'h103bc, 'h10973, 'h10974, 'h10975, 'h10976, 'h10001, 'h10000, 'h10977, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10978, 'h10979, 'h21f8c, 'h1097a, 'h1097b, 'h103bc, 'h1097c, 'h1097d, 'h1097e, 'h1097f, 'h10001, 'h10000, 'h10980, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10981, 'h10982, 'h21f8c, 'h10983, 'h10984, 'h103bc, 'h10985, 'h10986, 'h10987, 'h10988, 'h10001, 'h10000, 'h10989, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1098a, 'h1098b, 'h21f8c, 'h1098c, 'h1098d, 'h103bc, 'h1098e, 'h1098f, 'h10990, 'h10991, 'h10001, 'h10000, 'h10992, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10993, 'h10994, 'h21f8c, 'h10995, 'h10996, 'h103bc, 'h10997, 'h10998, 'h10999, 'h1099a, 'h10001, 'h10000, 'h1099b, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1099c, 'h1099d, 'h21f8c, 'h1099e, 'h1099f, 'h103bc, 'h109a0, 'h109a1, 'h109a2, 'h109a3, 'h10001, 'h10000, 'h109a4, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109a5, 'h109a6, 'h21f8c, 'h109a7, 'h109a8, 'h103bc, 'h109a9, 'h109aa, 'h109ab, 'h109ac, 'h10001, 'h10000, 'h109ad, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109ae, 'h109af, 'h21f8c, 'h109b0, 'h109b1, 'h103bc, 'h109b2, 'h109b3, 'h109b4, 'h109b5, 'h10001, 'h10000, 'h109b6, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109b7, 'h109b8, 'h21f8c, 'h109b9, 'h109ba, 'h103bc, 'h109bb, 'h109bc, 'h109bd, 'h109be, 'h10001, 'h10000, 'h109bf, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109c0, 'h109c1, 'h21f8c, 'h109c2, 'h109c3, 'h103bc, 'h109c4, 'h109c5, 'h109c6, 'h109c7, 'h10001, 'h10000, 'h109c8, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109c9, 'h109ca, 'h21f8c, 'h109cb, 'h109cc, 'h103bc, 'h109cd, 'h109ce, 'h109cf, 'h109d0, 'h10001, 'h10000, 'h109d1, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109d2, 'h109d3, 'h21f8c, 'h109d4, 'h109d5, 'h103bc, 'h109d6, 'h109d7, 'h109d8, 'h109d9, 'h10001, 'h10000, 'h109da, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109db, 'h109dc, 'h21f8c, 'h109dd, 'h109de, 'h103bc, 'h109df, 'h109e0, 'h109e1, 'h109e2, 'h10001, 'h10000, 'h109e3, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109e4, 'h109e5, 'h21f8c, 'h109e6, 'h109e7, 'h103bc, 'h109e8, 'h109e9, 'h109ea, 'h109eb, 'h10001, 'h10000, 'h109ec, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109ed, 'h109ee, 'h21f8c, 'h109ef, 'h109f0, 'h103bc, 'h109f1, 'h109f2, 'h109f3, 'h109f4, 'h10001, 'h10000, 'h109f5, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109f6, 'h109f7, 'h21f8c, 'h109f8, 'h109f9, 'h103bc, 'h109fa, 'h109fb, 'h109fc, 'h109fd, 'h10001, 'h10000, 'h109fe, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h109ff, 'h10a00, 'h21f8c, 'h10a01, 'h10a02, 'h103bc, 'h10a03, 'h10a04, 'h10a05, 'h10a06, 'h10001, 'h10000, 'h10a07, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a08, 'h10a09, 'h21f8c, 'h10a0a, 'h10a0b, 'h103bc, 'h10a0c, 'h10a0d, 'h10a0e, 'h10a0f, 'h10001, 'h10000, 'h10a10, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a11, 'h10a12, 'h21f8c, 'h10a13, 'h10a14, 'h103bc, 'h10a15, 'h10a16, 'h10a17, 'h10a18, 'h10001, 'h10000, 'h10a19, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a1a, 'h10a1b, 'h21f8c, 'h10a1c, 'h10a1d, 'h103bc, 'h10a1e, 'h10a1f, 'h10a20, 'h10a21, 'h10001, 'h10000, 'h10a22, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a23, 'h10a24, 'h21f8c, 'h10a25, 'h10a26, 'h103bc, 'h10a27, 'h10a28, 'h10a29, 'h10a2a, 'h10001, 'h10000, 'h10a2b, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a2c, 'h10a2d, 'h21f8c, 'h10a2e, 'h10a2f, 'h103bc, 'h10a30, 'h10a31, 'h10a32, 'h10a33, 'h10001, 'h10000, 'h10a34, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a35, 'h10a36, 'h21f8c, 'h10a37, 'h10a38, 'h103bc, 'h10a39, 'h10a3a, 'h10a3b, 'h10a3c, 'h10001, 'h10000, 'h10a3d, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a3e, 'h10a3f, 'h21f8c, 'h10a40, 'h10a41, 'h103bc, 'h10a42, 'h10a43, 'h10a44, 'h10a45, 'h10001, 'h10000, 'h10a46, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a47, 'h10a48, 'h21f8c, 'h10a49, 'h10a4a, 'h103bc, 'h10a4b, 'h10a4c, 'h10a4d, 'h10a4e, 'h10001, 'h10000, 'h10a4f, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a50, 'h10a51, 'h21f8c, 'h10a52, 'h10a53, 'h103bc, 'h10a54, 'h10a55, 'h10a56, 'h10a57, 'h10001, 'h10000, 'h10a58, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a59, 'h10a5a, 'h21f8c, 'h10a5b, 'h10a5c, 'h103bc, 'h10a5d, 'h10a5e, 'h10a5f, 'h10a60, 'h10001, 'h10000, 'h10a61, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a62, 'h10a63, 'h21f8c, 'h10a64, 'h10a65, 'h103bc, 'h10a66, 'h10a67, 'h10a68, 'h10a69, 'h10001, 'h10000, 'h10a6a, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a6b, 'h10a6c, 'h21f8c, 'h10a6d, 'h10a6e, 'h103bc, 'h10a6f, 'h10a70, 'h10a71, 'h10a72, 'h10001, 'h10000, 'h10a73, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a74, 'h10a75, 'h21f8c, 'h10a76, 'h10a77, 'h103bc, 'h10a78, 'h10a79, 'h10a7a, 'h10a7b, 'h10001, 'h10000, 'h10a7c, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a7d, 'h10a7e, 'h21f8c, 'h10a7f, 'h10a80, 'h103bc, 'h10a81, 'h10a82, 'h10a83, 'h10a84, 'h10001, 'h10000, 'h10a85, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a86, 'h10a87, 'h21f8c, 'h10a88, 'h10a89, 'h103bc, 'h10a8a, 'h10a8b, 'h10a8c, 'h10a8d, 'h10001, 'h10000, 'h10a8e, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a8f, 'h10a90, 'h21f8c, 'h10a91, 'h10a92, 'h103bc, 'h10a93, 'h10a94, 'h10a95, 'h10a96, 'h10001, 'h10000, 'h10a97, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10a98, 'h10a99, 'h21f8c, 'h10a9a, 'h10a9b, 'h103bc, 'h10a9c, 'h10a9d, 'h10a9e, 'h10a9f, 'h10001, 'h10000, 'h10aa0, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10aa1, 'h10aa2, 'h21f8c, 'h10aa3, 'h10aa4, 'h103bc, 'h10aa5, 'h10aa6, 'h10aa7, 'h10aa8, 'h10001, 'h10000, 'h10aa9, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10aaa, 'h10aab, 'h21f8c, 'h10aac, 'h10aad, 'h103bc, 'h10aae, 'h10aaf, 'h10ab0, 'h10ab1, 'h10001, 'h10000, 'h10ab2, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10ab3, 'h10ab4, 'h21f8c, 'h10ab5, 'h10ab6, 'h103bc, 'h10ab7, 'h10ab8, 'h10ab9, 'h10aba, 'h10001, 'h10000, 'h10abb, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10abc, 'h10abd, 'h21f8c, 'h10abe, 'h10abf, 'h103bc, 'h10ac0, 'h10ac1, 'h10ac2, 'h10ac3, 'h10001, 'h10000, 'h10ac4, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10ac5, 'h10ac6, 'h21f8c, 'h10ac7, 'h10ac8, 'h103bc, 'h10ac9, 'h10aca, 'h10acb, 'h10acc, 'h10001, 'h10000, 'h10acd, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10ace, 'h10acf, 'h21f8c, 'h10ad0, 'h10ad1, 'h103bc, 'h10ad2, 'h10ad3, 'h10ad4, 'h10ad5, 'h10001, 'h10000, 'h10ad6, 'h21f8b, 'h103bf, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10ad7, 'h10ad8, 'h21f8c, 'h10ad9, 'h10ada, 'h103bc, 'h10adb, 'h10adc, 'h10add, 'h21f8d, 'h10ade, 'h10adf, 'h10ae0, 'h21f8b, 'h10ae1, 'h10ae2, 'h10ae3, 'h10ae4, 'h10ae5, 'h10ae6, 'h10ae7, 'h10ae8, 'h10ae9, 'h10aea, 'h10aeb, 'h10aec, 'h103bc, 'h10aed, 'h10aee, 'h10aef, 'h10af0, 'h10af1, 'h10af2, 'h10af3, 'h21f8b, 'h10af4, 'h10af5, 'h10af6, 'h10af7, 'h10af8, 'h10af9, 'h10afa, 'h10afb, 'h10afc, 'h10afd, 'h10afe, 'h10aff, 'h103bc, 'h10b00, 'h10b01, 'h10b02, 'h10b03, 'h10b04, 'h10b05, 'h10b06, 'h21f8b, 'h10b07, 'h10b08, 'h10b09, 'h10b0a, 'h10b0b, 'h10b0c, 'h10b0d, 'h10b0e, 'h10b0f, 'h10b10, 'h10b11, 'h10b12, 'h103bc, 'h10b13, 'h10b14, 'h10b15, 'h10b16, 'h10b17, 'h10b18, 'h10b19, 'h21f8b, 'h10b1a, 'h10b1b, 'h10b1c, 'h10b1d, 'h10b1e, 'h10b1f, 'h10b20, 'h10b21, 'h10b22, 'h10b23, 'h10b24, 'h10b25, 'h103bc, 'h10b26, 'h10b27, 'h10b28, 'h10b29, 'h10b2a, 'h10b2b, 'h10b2c, 'h21f8b, 'h10b2d, 'h10b2e, 'h10b2f, 'h10b30, 'h10b31, 'h10b32, 'h10b33, 'h10b34, 'h10b35, 'h10b36, 'h10b37, 'h10b38, 'h103bc, 'h10b39, 'h10b3a, 'h10b3b, 'h10b3c, 'h10b3d, 'h10b3e, 'h10b3f, 'h21f8b, 'h10b40, 'h10b41, 'h10b42, 'h10b43, 'h10b44, 'h10b45, 'h10b46, 'h10b47, 'h10b48, 'h10b49, 'h10b4a, 'h10b4b, 'h103bc, 'h10b4c, 'h10b4d, 'h10b4e, 'h10b4f, 'h10b50, 'h10b51, 'h10b52, 'h21f8b, 'h10b53, 'h10b54, 'h10b55, 'h10b56, 'h10b57, 'h10b58, 'h10b59, 'h10b5a, 'h10b5b, 'h10b5c, 'h10b5d, 'h10b5e, 'h103bc, 'h10b5f, 'h10b60, 'h10b61, 'h10b62, 'h10b63, 'h10b64, 'h10b65, 'h21f8b, 'h10b66, 'h10b67, 'h10b68, 'h10b69, 'h10b6a, 'h10b6b, 'h10b6c, 'h10b6d, 'h10b6e, 'h10b6f, 'h10b70, 'h10b71, 'h103bc, 'h10b72, 'h10b73, 'h10b74, 'h10b75, 'h10b76, 'h10b77, 'h10b78, 'h21f8b, 'h10b79, 'h10b7a, 'h10b7b, 'h10b7c, 'h10b7d, 'h10b7e, 'h10b7f, 'h10b80, 'h10b81, 'h10b82, 'h10b83, 'h10b84, 'h103bc, 'h10b85, 'h10b86, 'h10b87, 'h10b88, 'h10b89, 'h10b8a, 'h10b8b, 'h21f8b, 'h10b8c, 'h10b8d, 'h10b8e, 'h10b8f, 'h10b90, 'h10b91, 'h10b92, 'h10b93, 'h10b94, 'h10b95, 'h10b96, 'h10b97, 'h103bc, 'h10b98, 'h10b99, 'h10b9a, 'h10b9b, 'h10b9c, 'h10b9d, 'h10b9e, 'h21f8b, 'h10b9f, 'h10ba0, 'h10ba1, 'h10ba2, 'h10ba3, 'h10ba4, 'h10ba5, 'h10ba6, 'h10ba7, 'h10ba8, 'h10ba9, 'h10baa, 'h103bc, 'h10bab, 'h10bac, 'h10bad, 'h10bae, 'h10baf, 'h10bb0, 'h10bb1, 'h21f8b, 'h10bb2, 'h10bb3, 'h10bb4, 'h10bb5, 'h10bb6, 'h10bb7, 'h10bb8, 'h10bb9, 'h10bba, 'h10bbb, 'h10bbc, 'h10bbd, 'h103bc, 'h10bbe, 'h10bbf, 'h10bc0, 'h10bc1, 'h10bc2, 'h10bc3, 'h10bc4, 'h21f8b, 'h10bc5, 'h10bc6, 'h10bc7, 'h10bc8, 'h10bc9, 'h10bca, 'h10bcb, 'h10bcc, 'h10bcd, 'h10bce, 'h10bcf, 'h10bd0, 'h103bc, 'h10bd1, 'h10bd2, 'h10bd3, 'h10bd4, 'h10bd5, 'h10bd6, 'h10bd7, 'h21f8b, 'h10bd8, 'h10bd9, 'h10bda, 'h10bdb, 'h10bdc, 'h10bdd, 'h10bde, 'h10bdf, 'h10be0, 'h10be1, 'h10be2, 'h10be3, 'h103bc, 'h10be4, 'h10be5, 'h10be6, 'h10be7, 'h10be8, 'h10be9, 'h10bea, 'h21f8b, 'h10beb, 'h10bec, 'h10bed, 'h10bee, 'h10bef, 'h10bf0, 'h10bf1, 'h10bf2, 'h10bf3, 'h10bf4, 'h10bf5, 'h10bf6, 'h103bc, 'h10bf7, 'h10bf8, 'h10bf9, 'h10bfa, 'h10bfb, 'h10bfc, 'h10bfd, 'h21f8b, 'h10bfe, 'h10bff, 'h10c00, 'h10c01, 'h10c02, 'h10c03, 'h10c04, 'h10c05, 'h10c06, 'h10c07, 'h10c08, 'h10c09, 'h103bc, 'h10c0a, 'h10c0b, 'h10c0c, 'h10c0d, 'h10c0e, 'h10c0f, 'h10c10, 'h21f8b, 'h10c11, 'h10c12, 'h10c13, 'h10c14, 'h10c15, 'h10c16, 'h10c17, 'h10c18, 'h10c19, 'h10c1a, 'h10c1b, 'h10c1c, 'h103bc, 'h10c1d, 'h10c1e, 'h10c1f, 'h10c20, 'h10c21, 'h10c22, 'h10c23, 'h21f8b, 'h10c24, 'h10c25, 'h10c26, 'h10c27, 'h10c28, 'h10c29, 'h10c2a, 'h10c2b, 'h10c2c, 'h10c2d, 'h10c2e, 'h10c2f, 'h103bc, 'h10c30, 'h10c31, 'h10c32, 'h10c33, 'h10c34, 'h10c35, 'h10c36, 'h21f8b, 'h10c37, 'h10c38, 'h10c39, 'h10c3a, 'h10c3b, 'h10c3c, 'h10c3d, 'h10c3e, 'h10c3f, 'h10c40, 'h10c41, 'h10c42, 'h103bc, 'h10c43, 'h10c44, 'h10c45, 'h10c46, 'h10c47, 'h10c48, 'h10c49, 'h21f8b, 'h10c4a, 'h10c4b, 'h10c4c, 'h10c4d, 'h10c4e, 'h10c4f, 'h10c50, 'h10c51, 'h10c52, 'h10c53, 'h10c54, 'h10c55, 'h103bc, 'h10c56, 'h10c57, 'h10c58, 'h10c59, 'h10c5a, 'h10c5b, 'h10c5c, 'h21f8b, 'h10c5d, 'h10c5e, 'h10c5f, 'h10c60, 'h10c61, 'h10c62, 'h10c63, 'h10c64, 'h10c65, 'h10c66, 'h10c67, 'h10c68, 'h103bc, 'h10c69, 'h10c6a, 'h10c6b, 'h10c6c, 'h10c6d, 'h10c6e, 'h10c6f, 'h21f8b, 'h10c70, 'h10c71, 'h10c72, 'h10c73, 'h10c74, 'h10c75, 'h10c76, 'h10c77, 'h10c78, 'h10c79, 'h10c7a, 'h10c7b, 'h103bc, 'h10c7c, 'h10c7d, 'h10c7e, 'h10c7f, 'h10c80, 'h10c81, 'h10c82, 'h21f8b, 'h10c83, 'h10c84, 'h10c85, 'h10c86, 'h10c87, 'h10c88, 'h10c89, 'h10c8a, 'h10c8b, 'h10c8c, 'h10c8d, 'h10c8e, 'h103bc, 'h10c8f, 'h10c90, 'h10c91, 'h10c92, 'h10c93, 'h10c94, 'h10c95, 'h21f8b, 'h10c96, 'h10c97, 'h10c98, 'h10c99, 'h10c9a, 'h10c9b, 'h10c9c, 'h10c9d, 'h10c9e, 'h10c9f, 'h10ca0, 'h10ca1, 'h103bc, 'h10ca2, 'h10ca3, 'h10ca4, 'h10ca5, 'h10ca6, 'h10ca7, 'h10ca8, 'h21f8b, 'h10ca9, 'h10caa, 'h10cab, 'h10cac, 'h10cad, 'h10cae, 'h10caf, 'h10cb0, 'h10cb1, 'h10cb2, 'h10cb3, 'h10cb4, 'h103bc, 'h10cb5, 'h10cb6, 'h10cb7, 'h10cb8, 'h10cb9, 'h10cba, 'h10cbb, 'h21f8b, 'h10cbc, 'h10cbd, 'h10cbe, 'h10cbf, 'h10cc0, 'h10cc1, 'h10cc2, 'h10cc3, 'h10cc4, 'h10cc5, 'h10cc6, 'h10cc7, 'h103bc, 'h10cc8, 'h10cc9, 'h10cca, 'h10ccb, 'h10ccc, 'h10ccd, 'h10cce, 'h21f8b, 'h10ccf, 'h10cd0, 'h10cd1, 'h10cd2, 'h10cd3, 'h10cd4, 'h10cd5, 'h10cd6, 'h10cd7, 'h10cd8, 'h10cd9, 'h10cda, 'h103bc, 'h10cdb, 'h10cdc, 'h10cdd, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h108de, 'h10ade, 'h106ee, 'h106fe, 'h108df, 'h1070e, 'h1071e, 'h108e0, 'h1072e, 'h1073e, 'h108e1, 'h1074e, 'h1075e, 'h108e2, 'h103bc, 'h1076e, 'h1077e, 'h108e3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078e, 'h10ade, 'h1079e, 'h108e4, 'h107ae, 'h107be, 'h108e5, 'h107ce, 'h107de, 'h108e6, 'h107ee, 'h107fe, 'h108e7, 'h1080e, 'h103bc, 'h1081e, 'h108e8, 'h1082e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083e, 'h108e9, 'h10ade, 'h1084e, 'h1085e, 'h108ea, 'h1086e, 'h1087e, 'h108eb, 'h1088e, 'h1089e, 'h108ec, 'h108ae, 'h108be, 'h108ed, 'h103bc, 'h108ce, 'h106de, 'h108ee, 'h10aee, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ee, 'h106fe, 'h108ef, 'h1070e, 'h1071e, 'h108f0, 'h1072e, 'h1073e, 'h108f1, 'h1074e, 'h1075e, 'h108f2, 'h1076e, 'h103bc, 'h1077e, 'h108f3, 'h1078e, 'h10aee, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079e, 'h108f4, 'h107ae, 'h107be, 'h108f5, 'h107ce, 'h107de, 'h108f6, 'h107ee, 'h107fe, 'h108f7, 'h1080e, 'h1081e, 'h108f8, 'h103bc, 'h1082e, 'h1083e, 'h108f9, 'h10aee, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084e, 'h1085e, 'h108fa, 'h1086e, 'h1087e, 'h108fb, 'h1088e, 'h1089e, 'h108fc, 'h108ae, 'h108be, 'h108fd, 'h108ce, 'h103bc, 'h106de, 'h108fe, 'h10afe, 'h106ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fe, 'h108ff, 'h1070e, 'h1071e, 'h10900, 'h1072e, 'h1073e, 'h10901, 'h1074e, 'h1075e, 'h10902, 'h1076e, 'h1077e, 'h10903, 'h103bc, 'h1078e, 'h10afe, 'h1079e, 'h10904, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ae, 'h107be, 'h10905, 'h107ce, 'h107de, 'h10906, 'h107ee, 'h107fe, 'h10907, 'h1080e, 'h1081e, 'h10908, 'h1082e, 'h103bc, 'h1083e, 'h10909, 'h10afe, 'h1084e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085e, 'h1090a, 'h1086e, 'h1087e, 'h1090b, 'h1088e, 'h1089e, 'h1090c, 'h108ae, 'h108be, 'h1090d, 'h108ce, 'h106de, 'h1090e, 'h10b0e, 'h103bc, 'h106ee, 'h106fe, 'h1090f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070e, 'h1071e, 'h10910, 'h1072e, 'h1073e, 'h10911, 'h1074e, 'h1075e, 'h10912, 'h1076e, 'h1077e, 'h10913, 'h1078e, 'h10b0e, 'h103bc, 'h1079e, 'h10914, 'h107ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h107be, 'h10915, 'h107ce, 'h107de, 'h10916, 'h107ee, 'h107fe, 'h10917, 'h1080e, 'h1081e, 'h10918, 'h1082e, 'h1083e, 'h10919, 'h10b0e, 'h103bc, 'h1084e, 'h1085e, 'h1091a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086e, 'h1087e, 'h1091b, 'h1088e, 'h1089e, 'h1091c, 'h108ae, 'h108be, 'h1091d, 'h108ce, 'h106de, 'h1091e, 'h10b1e, 'h106ee, 'h103bc, 'h106fe, 'h1091f, 'h1070e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071e, 'h10920, 'h1072e, 'h1073e, 'h10921, 'h1074e, 'h1075e, 'h10922, 'h1076e, 'h1077e, 'h10923, 'h1078e, 'h10b1e, 'h1079e, 'h10924, 'h103bc, 'h107ae, 'h107be, 'h10925, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ce, 'h107de, 'h10926, 'h107ee, 'h107fe, 'h10927, 'h1080e, 'h1081e, 'h10928, 'h1082e, 'h1083e, 'h10929, 'h10b1e, 'h1084e, 'h103bc, 'h1085e, 'h1092a, 'h1086e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087e, 'h1092b, 'h1088e, 'h1089e, 'h1092c, 'h108ae, 'h108be, 'h1092d, 'h108ce, 'h106de, 'h1092e, 'h10b2e, 'h106ee, 'h106fe, 'h1092f, 'h103bc, 'h1070e, 'h1071e, 'h10930, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072e, 'h1073e, 'h10931, 'h1074e, 'h1075e, 'h10932, 'h1076e, 'h1077e, 'h10933, 'h1078e, 'h10b2e, 'h1079e, 'h10934, 'h107ae, 'h103bc, 'h107be, 'h10935, 'h107ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h107de, 'h10936, 'h107ee, 'h107fe, 'h10937, 'h1080e, 'h1081e, 'h10938, 'h1082e, 'h1083e, 'h10939, 'h10b2e, 'h1084e, 'h1085e, 'h1093a, 'h103bc, 'h1086e, 'h1087e, 'h1093b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088e, 'h1089e, 'h1093c, 'h108ae, 'h108be, 'h1093d, 'h108ce, 'h106de, 'h1093e, 'h10b3e, 'h106ee, 'h106fe, 'h1093f, 'h1070e, 'h103bc, 'h1071e, 'h10940, 'h1072e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073e, 'h10941, 'h1074e, 'h1075e, 'h10942, 'h1076e, 'h1077e, 'h10943, 'h1078e, 'h10b3e, 'h1079e, 'h10944, 'h107ae, 'h107be, 'h10945, 'h103bc, 'h107ce, 'h107de, 'h10946, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ee, 'h107fe, 'h10947, 'h1080e, 'h1081e, 'h10948, 'h1082e, 'h1083e, 'h10949, 'h10b3e, 'h1084e, 'h1085e, 'h1094a, 'h1086e, 'h103bc, 'h1087e, 'h1094b, 'h1088e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089e, 'h1094c, 'h108ae, 'h108be, 'h1094d, 'h108ce, 'h106de, 'h1094e, 'h10b4e, 'h106ee, 'h106fe, 'h1094f, 'h1070e, 'h1071e, 'h10950, 'h103bc, 'h1072e, 'h1073e, 'h10951, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074e, 'h1075e, 'h10952, 'h1076e, 'h1077e, 'h10953, 'h1078e, 'h10b4e, 'h1079e, 'h10954, 'h107ae, 'h107be, 'h10955, 'h107ce, 'h103bc, 'h107de, 'h10956, 'h107ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fe, 'h10957, 'h1080e, 'h1081e, 'h10958, 'h1082e, 'h1083e, 'h10959, 'h10b4e, 'h1084e, 'h1085e, 'h1095a, 'h1086e, 'h1087e, 'h1095b, 'h103bc, 'h1088e, 'h1089e, 'h1095c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ae, 'h108be, 'h1095d, 'h108ce, 'h106de, 'h1095e, 'h10b5e, 'h106ee, 'h106fe, 'h1095f, 'h1070e, 'h1071e, 'h10960, 'h1072e, 'h103bc, 'h1073e, 'h10961, 'h1074e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075e, 'h10962, 'h1076e, 'h1077e, 'h10963, 'h1078e, 'h10b5e, 'h1079e, 'h10964, 'h107ae, 'h107be, 'h10965, 'h107ce, 'h107de, 'h10966, 'h103bc, 'h107ee, 'h107fe, 'h10967, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080e, 'h1081e, 'h10968, 'h1082e, 'h1083e, 'h10969, 'h10b5e, 'h1084e, 'h1085e, 'h1096a, 'h1086e, 'h1087e, 'h1096b, 'h1088e, 'h103bc, 'h1089e, 'h1096c, 'h108ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h108be, 'h1096d, 'h108ce, 'h106de, 'h1096e, 'h10b6e, 'h106ee, 'h106fe, 'h1096f, 'h1070e, 'h1071e, 'h10970, 'h1072e, 'h1073e, 'h10971, 'h103bc, 'h1074e, 'h1075e, 'h10972, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076e, 'h1077e, 'h10973, 'h1078e, 'h10b6e, 'h1079e, 'h10974, 'h107ae, 'h107be, 'h10975, 'h107ce, 'h107de, 'h10976, 'h107ee, 'h103bc, 'h107fe, 'h10977, 'h1080e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081e, 'h10978, 'h1082e, 'h1083e, 'h10979, 'h10b6e, 'h1084e, 'h1085e, 'h1097a, 'h1086e, 'h1087e, 'h1097b, 'h1088e, 'h1089e, 'h1097c, 'h103bc, 'h108ae, 'h108be, 'h1097d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ce, 'h106de, 'h1097e, 'h10b7e, 'h106ee, 'h106fe, 'h1097f, 'h1070e, 'h1071e, 'h10980, 'h1072e, 'h1073e, 'h10981, 'h1074e, 'h103bc, 'h1075e, 'h10982, 'h1076e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077e, 'h10983, 'h1078e, 'h10b7e, 'h1079e, 'h10984, 'h107ae, 'h107be, 'h10985, 'h107ce, 'h107de, 'h10986, 'h107ee, 'h107fe, 'h10987, 'h103bc, 'h1080e, 'h1081e, 'h10988, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082e, 'h1083e, 'h10989, 'h10b7e, 'h1084e, 'h1085e, 'h1098a, 'h1086e, 'h1087e, 'h1098b, 'h1088e, 'h1089e, 'h1098c, 'h108ae, 'h103bc, 'h108be, 'h1098d, 'h108ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1098e, 'h10b8e, 'h106ee, 'h106fe, 'h1098f, 'h1070e, 'h1071e, 'h10990, 'h1072e, 'h1073e, 'h10991, 'h1074e, 'h1075e, 'h10992, 'h103bc, 'h1076e, 'h1077e, 'h10993, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078e, 'h10b8e, 'h1079e, 'h10994, 'h107ae, 'h107be, 'h10995, 'h107ce, 'h107de, 'h10996, 'h107ee, 'h107fe, 'h10997, 'h1080e, 'h103bc, 'h1081e, 'h10998, 'h1082e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083e, 'h10999, 'h10b8e, 'h1084e, 'h1085e, 'h1099a, 'h1086e, 'h1087e, 'h1099b, 'h1088e, 'h1089e, 'h1099c, 'h108ae, 'h108be, 'h1099d, 'h103bc, 'h108ce, 'h106de, 'h1099e, 'h10b9e, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ee, 'h106fe, 'h1099f, 'h1070e, 'h1071e, 'h109a0, 'h1072e, 'h1073e, 'h109a1, 'h1074e, 'h1075e, 'h109a2, 'h1076e, 'h103bc, 'h1077e, 'h109a3, 'h1078e, 'h10b9e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079e, 'h109a4, 'h107ae, 'h107be, 'h109a5, 'h107ce, 'h107de, 'h109a6, 'h107ee, 'h107fe, 'h109a7, 'h1080e, 'h1081e, 'h109a8, 'h103bc, 'h1082e, 'h1083e, 'h109a9, 'h10b9e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084e, 'h1085e, 'h109aa, 'h1086e, 'h1087e, 'h109ab, 'h1088e, 'h1089e, 'h109ac, 'h108ae, 'h108be, 'h109ad, 'h108ce, 'h103bc, 'h106de, 'h109ae, 'h10bae, 'h106ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fe, 'h109af, 'h1070e, 'h1071e, 'h109b0, 'h1072e, 'h1073e, 'h109b1, 'h1074e, 'h1075e, 'h109b2, 'h1076e, 'h1077e, 'h109b3, 'h103bc, 'h1078e, 'h10bae, 'h1079e, 'h109b4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ae, 'h107be, 'h109b5, 'h107ce, 'h107de, 'h109b6, 'h107ee, 'h107fe, 'h109b7, 'h1080e, 'h1081e, 'h109b8, 'h1082e, 'h103bc, 'h1083e, 'h109b9, 'h10bae, 'h1084e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085e, 'h109ba, 'h1086e, 'h1087e, 'h109bb, 'h1088e, 'h1089e, 'h109bc, 'h108ae, 'h108be, 'h109bd, 'h108ce, 'h106de, 'h109be, 'h10bbe, 'h103bc, 'h106ee, 'h106fe, 'h109bf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070e, 'h1071e, 'h109c0, 'h1072e, 'h1073e, 'h109c1, 'h1074e, 'h1075e, 'h109c2, 'h1076e, 'h1077e, 'h109c3, 'h1078e, 'h10bbe, 'h103bc, 'h1079e, 'h109c4, 'h107ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h107be, 'h109c5, 'h107ce, 'h107de, 'h109c6, 'h107ee, 'h107fe, 'h109c7, 'h1080e, 'h1081e, 'h109c8, 'h1082e, 'h1083e, 'h109c9, 'h10bbe, 'h103bc, 'h1084e, 'h1085e, 'h109ca, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086e, 'h1087e, 'h109cb, 'h1088e, 'h1089e, 'h109cc, 'h108ae, 'h108be, 'h109cd, 'h108ce, 'h106de, 'h109ce, 'h10bce, 'h106ee, 'h103bc, 'h106fe, 'h109cf, 'h1070e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071e, 'h109d0, 'h1072e, 'h1073e, 'h109d1, 'h1074e, 'h1075e, 'h109d2, 'h1076e, 'h1077e, 'h109d3, 'h1078e, 'h10bce, 'h1079e, 'h109d4, 'h103bc, 'h107ae, 'h107be, 'h109d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ce, 'h107de, 'h109d6, 'h107ee, 'h107fe, 'h109d7, 'h1080e, 'h1081e, 'h109d8, 'h1082e, 'h1083e, 'h109d9, 'h10bce, 'h1084e, 'h103bc, 'h1085e, 'h109da, 'h1086e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087e, 'h109db, 'h1088e, 'h1089e, 'h109dc, 'h108ae, 'h108be, 'h109dd, 'h108ce, 'h106de, 'h109de, 'h10bde, 'h106ee, 'h106fe, 'h109df, 'h103bc, 'h1070e, 'h1071e, 'h109e0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072e, 'h1073e, 'h109e1, 'h1074e, 'h1075e, 'h109e2, 'h1076e, 'h1077e, 'h109e3, 'h1078e, 'h10bde, 'h1079e, 'h109e4, 'h107ae, 'h103bc, 'h107be, 'h109e5, 'h107ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h107de, 'h109e6, 'h107ee, 'h107fe, 'h109e7, 'h1080e, 'h1081e, 'h109e8, 'h1082e, 'h1083e, 'h109e9, 'h10bde, 'h1084e, 'h1085e, 'h109ea, 'h103bc, 'h1086e, 'h1087e, 'h109eb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088e, 'h1089e, 'h109ec, 'h108ae, 'h108be, 'h109ed, 'h108ce, 'h106de, 'h109ee, 'h10bee, 'h106ee, 'h106fe, 'h109ef, 'h1070e, 'h103bc, 'h1071e, 'h109f0, 'h1072e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073e, 'h109f1, 'h1074e, 'h1075e, 'h109f2, 'h1076e, 'h1077e, 'h109f3, 'h1078e, 'h10bee, 'h1079e, 'h109f4, 'h107ae, 'h107be, 'h109f5, 'h103bc, 'h107ce, 'h107de, 'h109f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ee, 'h107fe, 'h109f7, 'h1080e, 'h1081e, 'h109f8, 'h1082e, 'h1083e, 'h109f9, 'h10bee, 'h1084e, 'h1085e, 'h109fa, 'h1086e, 'h103bc, 'h1087e, 'h109fb, 'h1088e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089e, 'h109fc, 'h108ae, 'h108be, 'h109fd, 'h108ce, 'h106de, 'h109fe, 'h10bfe, 'h106ee, 'h106fe, 'h109ff, 'h1070e, 'h1071e, 'h10a00, 'h103bc, 'h1072e, 'h1073e, 'h10a01, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074e, 'h1075e, 'h10a02, 'h1076e, 'h1077e, 'h10a03, 'h1078e, 'h10bfe, 'h1079e, 'h10a04, 'h107ae, 'h107be, 'h10a05, 'h107ce, 'h103bc, 'h107de, 'h10a06, 'h107ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fe, 'h10a07, 'h1080e, 'h1081e, 'h10a08, 'h1082e, 'h1083e, 'h10a09, 'h10bfe, 'h1084e, 'h1085e, 'h10a0a, 'h1086e, 'h1087e, 'h10a0b, 'h103bc, 'h1088e, 'h1089e, 'h10a0c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ae, 'h108be, 'h10a0d, 'h108ce, 'h106de, 'h10a0e, 'h10c0e, 'h106ee, 'h106fe, 'h10a0f, 'h1070e, 'h1071e, 'h10a10, 'h1072e, 'h103bc, 'h1073e, 'h10a11, 'h1074e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075e, 'h10a12, 'h1076e, 'h1077e, 'h10a13, 'h1078e, 'h10c0e, 'h1079e, 'h10a14, 'h107ae, 'h107be, 'h10a15, 'h107ce, 'h107de, 'h10a16, 'h103bc, 'h107ee, 'h107fe, 'h10a17, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080e, 'h1081e, 'h10a18, 'h1082e, 'h1083e, 'h10a19, 'h10c0e, 'h1084e, 'h1085e, 'h10a1a, 'h1086e, 'h1087e, 'h10a1b, 'h1088e, 'h103bc, 'h1089e, 'h10a1c, 'h108ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h108be, 'h10a1d, 'h108ce, 'h106de, 'h10a1e, 'h10c1e, 'h106ee, 'h106fe, 'h10a1f, 'h1070e, 'h1071e, 'h10a20, 'h1072e, 'h1073e, 'h10a21, 'h103bc, 'h1074e, 'h1075e, 'h10a22, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076e, 'h1077e, 'h10a23, 'h1078e, 'h10c1e, 'h1079e, 'h10a24, 'h107ae, 'h107be, 'h10a25, 'h107ce, 'h107de, 'h10a26, 'h107ee, 'h103bc, 'h107fe, 'h10a27, 'h1080e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081e, 'h10a28, 'h1082e, 'h1083e, 'h10a29, 'h10c1e, 'h1084e, 'h1085e, 'h10a2a, 'h1086e, 'h1087e, 'h10a2b, 'h1088e, 'h1089e, 'h10a2c, 'h103bc, 'h108ae, 'h108be, 'h10a2d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ce, 'h106de, 'h10a2e, 'h10c2e, 'h106ee, 'h106fe, 'h10a2f, 'h1070e, 'h1071e, 'h10a30, 'h1072e, 'h1073e, 'h10a31, 'h1074e, 'h103bc, 'h1075e, 'h10a32, 'h1076e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077e, 'h10a33, 'h1078e, 'h10c2e, 'h1079e, 'h10a34, 'h107ae, 'h107be, 'h10a35, 'h107ce, 'h107de, 'h10a36, 'h107ee, 'h107fe, 'h10a37, 'h103bc, 'h1080e, 'h1081e, 'h10a38, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082e, 'h1083e, 'h10a39, 'h10c2e, 'h1084e, 'h1085e, 'h10a3a, 'h1086e, 'h1087e, 'h10a3b, 'h1088e, 'h1089e, 'h10a3c, 'h108ae, 'h103bc, 'h108be, 'h10a3d, 'h108ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h10a3e, 'h10c3e, 'h106ee, 'h106fe, 'h10a3f, 'h1070e, 'h1071e, 'h10a40, 'h1072e, 'h1073e, 'h10a41, 'h1074e, 'h1075e, 'h10a42, 'h103bc, 'h1076e, 'h1077e, 'h10a43, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078e, 'h10c3e, 'h1079e, 'h10a44, 'h107ae, 'h107be, 'h10a45, 'h107ce, 'h107de, 'h10a46, 'h107ee, 'h107fe, 'h10a47, 'h1080e, 'h103bc, 'h1081e, 'h10a48, 'h1082e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083e, 'h10a49, 'h10c3e, 'h1084e, 'h1085e, 'h10a4a, 'h1086e, 'h1087e, 'h10a4b, 'h1088e, 'h1089e, 'h10a4c, 'h108ae, 'h108be, 'h10a4d, 'h103bc, 'h108ce, 'h106de, 'h10a4e, 'h10c4e, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ee, 'h106fe, 'h10a4f, 'h1070e, 'h1071e, 'h10a50, 'h1072e, 'h1073e, 'h10a51, 'h1074e, 'h1075e, 'h10a52, 'h1076e, 'h103bc, 'h1077e, 'h10a53, 'h1078e, 'h10c4e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079e, 'h10a54, 'h107ae, 'h107be, 'h10a55, 'h107ce, 'h107de, 'h10a56, 'h107ee, 'h107fe, 'h10a57, 'h1080e, 'h1081e, 'h10a58, 'h103bc, 'h1082e, 'h1083e, 'h10a59, 'h10c4e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084e, 'h1085e, 'h10a5a, 'h1086e, 'h1087e, 'h10a5b, 'h1088e, 'h1089e, 'h10a5c, 'h108ae, 'h108be, 'h10a5d, 'h108ce, 'h103bc, 'h106de, 'h10a5e, 'h10c5e, 'h106ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fe, 'h10a5f, 'h1070e, 'h1071e, 'h10a60, 'h1072e, 'h1073e, 'h10a61, 'h1074e, 'h1075e, 'h10a62, 'h1076e, 'h1077e, 'h10a63, 'h103bc, 'h1078e, 'h10c5e, 'h1079e, 'h10a64, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ae, 'h107be, 'h10a65, 'h107ce, 'h107de, 'h10a66, 'h107ee, 'h107fe, 'h10a67, 'h1080e, 'h1081e, 'h10a68, 'h1082e, 'h103bc, 'h1083e, 'h10a69, 'h10c5e, 'h1084e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085e, 'h10a6a, 'h1086e, 'h1087e, 'h10a6b, 'h1088e, 'h1089e, 'h10a6c, 'h108ae, 'h108be, 'h10a6d, 'h108ce, 'h106de, 'h10a6e, 'h10c6e, 'h103bc, 'h106ee, 'h106fe, 'h10a6f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070e, 'h1071e, 'h10a70, 'h1072e, 'h1073e, 'h10a71, 'h1074e, 'h1075e, 'h10a72, 'h1076e, 'h1077e, 'h10a73, 'h1078e, 'h10c6e, 'h103bc, 'h1079e, 'h10a74, 'h107ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h107be, 'h10a75, 'h107ce, 'h107de, 'h10a76, 'h107ee, 'h107fe, 'h10a77, 'h1080e, 'h1081e, 'h10a78, 'h1082e, 'h1083e, 'h10a79, 'h10c6e, 'h103bc, 'h1084e, 'h1085e, 'h10a7a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086e, 'h1087e, 'h10a7b, 'h1088e, 'h1089e, 'h10a7c, 'h108ae, 'h108be, 'h10a7d, 'h108ce, 'h106de, 'h10a7e, 'h10c7e, 'h106ee, 'h103bc, 'h106fe, 'h10a7f, 'h1070e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071e, 'h10a80, 'h1072e, 'h1073e, 'h10a81, 'h1074e, 'h1075e, 'h10a82, 'h1076e, 'h1077e, 'h10a83, 'h1078e, 'h10c7e, 'h1079e, 'h10a84, 'h103bc, 'h107ae, 'h107be, 'h10a85, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ce, 'h107de, 'h10a86, 'h107ee, 'h107fe, 'h10a87, 'h1080e, 'h1081e, 'h10a88, 'h1082e, 'h1083e, 'h10a89, 'h10c7e, 'h1084e, 'h103bc, 'h1085e, 'h10a8a, 'h1086e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087e, 'h10a8b, 'h1088e, 'h1089e, 'h10a8c, 'h108ae, 'h108be, 'h10a8d, 'h108ce, 'h106de, 'h10a8e, 'h10c8e, 'h106ee, 'h106fe, 'h10a8f, 'h103bc, 'h1070e, 'h1071e, 'h10a90, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072e, 'h1073e, 'h10a91, 'h1074e, 'h1075e, 'h10a92, 'h1076e, 'h1077e, 'h10a93, 'h1078e, 'h10c8e, 'h1079e, 'h10a94, 'h107ae, 'h103bc, 'h107be, 'h10a95, 'h107ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h107de, 'h10a96, 'h107ee, 'h107fe, 'h10a97, 'h1080e, 'h1081e, 'h10a98, 'h1082e, 'h1083e, 'h10a99, 'h10c8e, 'h1084e, 'h1085e, 'h10a9a, 'h103bc, 'h1086e, 'h1087e, 'h10a9b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088e, 'h1089e, 'h10a9c, 'h108ae, 'h108be, 'h10a9d, 'h108ce, 'h106de, 'h10a9e, 'h10c9e, 'h106ee, 'h106fe, 'h10a9f, 'h1070e, 'h103bc, 'h1071e, 'h10aa0, 'h1072e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073e, 'h10aa1, 'h1074e, 'h1075e, 'h10aa2, 'h1076e, 'h1077e, 'h10aa3, 'h1078e, 'h10c9e, 'h1079e, 'h10aa4, 'h107ae, 'h107be, 'h10aa5, 'h103bc, 'h107ce, 'h107de, 'h10aa6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ee, 'h107fe, 'h10aa7, 'h1080e, 'h1081e, 'h10aa8, 'h1082e, 'h1083e, 'h10aa9, 'h10c9e, 'h1084e, 'h1085e, 'h10aaa, 'h1086e, 'h103bc, 'h1087e, 'h10aab, 'h1088e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089e, 'h10aac, 'h108ae, 'h108be, 'h10aad, 'h108ce, 'h106de, 'h10aae, 'h10cae, 'h106ee, 'h106fe, 'h10aaf, 'h1070e, 'h1071e, 'h10ab0, 'h103bc, 'h1072e, 'h1073e, 'h10ab1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074e, 'h1075e, 'h10ab2, 'h1076e, 'h1077e, 'h10ab3, 'h1078e, 'h10cae, 'h1079e, 'h10ab4, 'h107ae, 'h107be, 'h10ab5, 'h107ce, 'h103bc, 'h107de, 'h10ab6, 'h107ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fe, 'h10ab7, 'h1080e, 'h1081e, 'h10ab8, 'h1082e, 'h1083e, 'h10ab9, 'h10cae, 'h1084e, 'h1085e, 'h10aba, 'h1086e, 'h1087e, 'h10abb, 'h103bc, 'h1088e, 'h1089e, 'h10abc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ae, 'h108be, 'h10abd, 'h108ce, 'h106de, 'h10abe, 'h10cbe, 'h106ee, 'h106fe, 'h10abf, 'h1070e, 'h1071e, 'h10ac0, 'h1072e, 'h103bc, 'h1073e, 'h10ac1, 'h1074e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075e, 'h10ac2, 'h1076e, 'h1077e, 'h10ac3, 'h1078e, 'h10cbe, 'h1079e, 'h10ac4, 'h107ae, 'h107be, 'h10ac5, 'h107ce, 'h107de, 'h10ac6, 'h103bc, 'h107ee, 'h107fe, 'h10ac7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080e, 'h1081e, 'h10ac8, 'h1082e, 'h1083e, 'h10ac9, 'h10cbe, 'h1084e, 'h1085e, 'h10aca, 'h1086e, 'h1087e, 'h10acb, 'h1088e, 'h103bc, 'h1089e, 'h10acc, 'h108ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h108be, 'h10acd, 'h108ce, 'h106de, 'h10ace, 'h10cce, 'h106ee, 'h106fe, 'h10acf, 'h1070e, 'h1071e, 'h10ad0, 'h1072e, 'h1073e, 'h10ad1, 'h103bc, 'h1074e, 'h1075e, 'h10ad2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076e, 'h1077e, 'h10ad3, 'h1078e, 'h10cce, 'h1079e, 'h10ad4, 'h107ae, 'h107be, 'h10ad5, 'h107ce, 'h107de, 'h10ad6, 'h107ee, 'h103bc, 'h107fe, 'h10ad7, 'h1080e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081e, 'h10ad8, 'h1082e, 'h1083e, 'h10ad9, 'h10cce, 'h1084e, 'h1085e, 'h10ada, 'h1086e, 'h1087e, 'h10adb, 'h1088e, 'h1089e, 'h10adc, 'h103bc, 'h108ae, 'h108be, 'h10add, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ce, 'h106de, 'h108de, 'h10ade, 'h106ee, 'h106fe, 'h108df, 'h1070e, 'h1071e, 'h108e0, 'h1072e, 'h1073e, 'h108e1, 'h1074e, 'h103bc, 'h1075e, 'h108e2, 'h1076e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077e, 'h108e3, 'h1078e, 'h10ade, 'h1079e, 'h108e4, 'h107ae, 'h107be, 'h108e5, 'h107ce, 'h107de, 'h108e6, 'h107ee, 'h107fe, 'h108e7, 'h103bc, 'h1080e, 'h1081e, 'h108e8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082e, 'h1083e, 'h108e9, 'h10ade, 'h1084e, 'h1085e, 'h108ea, 'h1086e, 'h1087e, 'h108eb, 'h1088e, 'h1089e, 'h108ec, 'h108ae, 'h103bc, 'h108be, 'h108ed, 'h108ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h108ee, 'h10aee, 'h106ee, 'h106fe, 'h108ef, 'h1070e, 'h1071e, 'h108f0, 'h1072e, 'h1073e, 'h108f1, 'h1074e, 'h1075e, 'h108f2, 'h103bc, 'h1076e, 'h1077e, 'h108f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078e, 'h10aee, 'h1079e, 'h108f4, 'h107ae, 'h107be, 'h108f5, 'h107ce, 'h107de, 'h108f6, 'h107ee, 'h107fe, 'h108f7, 'h1080e, 'h103bc, 'h1081e, 'h108f8, 'h1082e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083e, 'h108f9, 'h10aee, 'h1084e, 'h1085e, 'h108fa, 'h1086e, 'h1087e, 'h108fb, 'h1088e, 'h1089e, 'h108fc, 'h108ae, 'h108be, 'h108fd, 'h103bc, 'h108ce, 'h106de, 'h108fe, 'h10afe, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ee, 'h106fe, 'h108ff, 'h1070e, 'h1071e, 'h10900, 'h1072e, 'h1073e, 'h10901, 'h1074e, 'h1075e, 'h10902, 'h1076e, 'h103bc, 'h1077e, 'h10903, 'h1078e, 'h10afe, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079e, 'h10904, 'h107ae, 'h107be, 'h10905, 'h107ce, 'h107de, 'h10906, 'h107ee, 'h107fe, 'h10907, 'h1080e, 'h1081e, 'h10908, 'h103bc, 'h1082e, 'h1083e, 'h10909, 'h10afe, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084e, 'h1085e, 'h1090a, 'h1086e, 'h1087e, 'h1090b, 'h1088e, 'h1089e, 'h1090c, 'h108ae, 'h108be, 'h1090d, 'h108ce, 'h103bc, 'h106de, 'h1090e, 'h10b0e, 'h106ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fe, 'h1090f, 'h1070e, 'h1071e, 'h10910, 'h1072e, 'h1073e, 'h10911, 'h1074e, 'h1075e, 'h10912, 'h1076e, 'h1077e, 'h10913, 'h103bc, 'h1078e, 'h10b0e, 'h1079e, 'h10914, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ae, 'h107be, 'h10915, 'h107ce, 'h107de, 'h10916, 'h107ee, 'h107fe, 'h10917, 'h1080e, 'h1081e, 'h10918, 'h1082e, 'h103bc, 'h1083e, 'h10919, 'h10b0e, 'h1084e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085e, 'h1091a, 'h1086e, 'h1087e, 'h1091b, 'h1088e, 'h1089e, 'h1091c, 'h108ae, 'h108be, 'h1091d, 'h108ce, 'h106de, 'h1091e, 'h10b1e, 'h103bc, 'h106ee, 'h106fe, 'h1091f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070e, 'h1071e, 'h10920, 'h1072e, 'h1073e, 'h10921, 'h1074e, 'h1075e, 'h10922, 'h1076e, 'h1077e, 'h10923, 'h1078e, 'h10b1e, 'h103bc, 'h1079e, 'h10924, 'h107ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h107be, 'h10925, 'h107ce, 'h107de, 'h10926, 'h107ee, 'h107fe, 'h10927, 'h1080e, 'h1081e, 'h10928, 'h1082e, 'h1083e, 'h10929, 'h10b1e, 'h103bc, 'h1084e, 'h1085e, 'h1092a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086e, 'h1087e, 'h1092b, 'h1088e, 'h1089e, 'h1092c, 'h108ae, 'h108be, 'h1092d, 'h108ce, 'h106de, 'h1092e, 'h10b2e, 'h106ee, 'h103bc, 'h106fe, 'h1092f, 'h1070e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071e, 'h10930, 'h1072e, 'h1073e, 'h10931, 'h1074e, 'h1075e, 'h10932, 'h1076e, 'h1077e, 'h10933, 'h1078e, 'h10b2e, 'h1079e, 'h10934, 'h103bc, 'h107ae, 'h107be, 'h10935, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ce, 'h107de, 'h10936, 'h107ee, 'h107fe, 'h10937, 'h1080e, 'h1081e, 'h10938, 'h1082e, 'h1083e, 'h10939, 'h10b2e, 'h1084e, 'h103bc, 'h1085e, 'h1093a, 'h1086e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087e, 'h1093b, 'h1088e, 'h1089e, 'h1093c, 'h108ae, 'h108be, 'h1093d, 'h108ce, 'h106de, 'h1093e, 'h10b3e, 'h106ee, 'h106fe, 'h1093f, 'h103bc, 'h1070e, 'h1071e, 'h10940, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072e, 'h1073e, 'h10941, 'h1074e, 'h1075e, 'h10942, 'h1076e, 'h1077e, 'h10943, 'h1078e, 'h10b3e, 'h1079e, 'h10944, 'h107ae, 'h103bc, 'h107be, 'h10945, 'h107ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h107de, 'h10946, 'h107ee, 'h107fe, 'h10947, 'h1080e, 'h1081e, 'h10948, 'h1082e, 'h1083e, 'h10949, 'h10b3e, 'h1084e, 'h1085e, 'h1094a, 'h103bc, 'h1086e, 'h1087e, 'h1094b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088e, 'h1089e, 'h1094c, 'h108ae, 'h108be, 'h1094d, 'h108ce, 'h106de, 'h1094e, 'h10b4e, 'h106ee, 'h106fe, 'h1094f, 'h1070e, 'h103bc, 'h1071e, 'h10950, 'h1072e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073e, 'h10951, 'h1074e, 'h1075e, 'h10952, 'h1076e, 'h1077e, 'h10953, 'h1078e, 'h10b4e, 'h1079e, 'h10954, 'h107ae, 'h107be, 'h10955, 'h103bc, 'h107ce, 'h107de, 'h10956, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ee, 'h107fe, 'h10957, 'h1080e, 'h1081e, 'h10958, 'h1082e, 'h1083e, 'h10959, 'h10b4e, 'h1084e, 'h1085e, 'h1095a, 'h1086e, 'h103bc, 'h1087e, 'h1095b, 'h1088e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089e, 'h1095c, 'h108ae, 'h108be, 'h1095d, 'h108ce, 'h106de, 'h1095e, 'h10b5e, 'h106ee, 'h106fe, 'h1095f, 'h1070e, 'h1071e, 'h10960, 'h103bc, 'h1072e, 'h1073e, 'h10961, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074e, 'h1075e, 'h10962, 'h1076e, 'h1077e, 'h10963, 'h1078e, 'h10b5e, 'h1079e, 'h10964, 'h107ae, 'h107be, 'h10965, 'h107ce, 'h103bc, 'h107de, 'h10966, 'h107ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fe, 'h10967, 'h1080e, 'h1081e, 'h10968, 'h1082e, 'h1083e, 'h10969, 'h10b5e, 'h1084e, 'h1085e, 'h1096a, 'h1086e, 'h1087e, 'h1096b, 'h103bc, 'h1088e, 'h1089e, 'h1096c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ae, 'h108be, 'h1096d, 'h108ce, 'h106de, 'h1096e, 'h10b6e, 'h106ee, 'h106fe, 'h1096f, 'h1070e, 'h1071e, 'h10970, 'h1072e, 'h103bc, 'h1073e, 'h10971, 'h1074e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075e, 'h10972, 'h1076e, 'h1077e, 'h10973, 'h1078e, 'h10b6e, 'h1079e, 'h10974, 'h107ae, 'h107be, 'h10975, 'h107ce, 'h107de, 'h10976, 'h103bc, 'h107ee, 'h107fe, 'h10977, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080e, 'h1081e, 'h10978, 'h1082e, 'h1083e, 'h10979, 'h10b6e, 'h1084e, 'h1085e, 'h1097a, 'h1086e, 'h1087e, 'h1097b, 'h1088e, 'h103bc, 'h1089e, 'h1097c, 'h108ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h108be, 'h1097d, 'h108ce, 'h106de, 'h1097e, 'h10b7e, 'h106ee, 'h106fe, 'h1097f, 'h1070e, 'h1071e, 'h10980, 'h1072e, 'h1073e, 'h10981, 'h103bc, 'h1074e, 'h1075e, 'h10982, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076e, 'h1077e, 'h10983, 'h1078e, 'h10b7e, 'h1079e, 'h10984, 'h107ae, 'h107be, 'h10985, 'h107ce, 'h107de, 'h10986, 'h107ee, 'h103bc, 'h107fe, 'h10987, 'h1080e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081e, 'h10988, 'h1082e, 'h1083e, 'h10989, 'h10b7e, 'h1084e, 'h1085e, 'h1098a, 'h1086e, 'h1087e, 'h1098b, 'h1088e, 'h1089e, 'h1098c, 'h103bc, 'h108ae, 'h108be, 'h1098d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ce, 'h106de, 'h1098e, 'h10b8e, 'h106ee, 'h106fe, 'h1098f, 'h1070e, 'h1071e, 'h10990, 'h1072e, 'h1073e, 'h10991, 'h1074e, 'h103bc, 'h1075e, 'h10992, 'h1076e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077e, 'h10993, 'h1078e, 'h10b8e, 'h1079e, 'h10994, 'h107ae, 'h107be, 'h10995, 'h107ce, 'h107de, 'h10996, 'h107ee, 'h107fe, 'h10997, 'h103bc, 'h1080e, 'h1081e, 'h10998, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082e, 'h1083e, 'h10999, 'h10b8e, 'h1084e, 'h1085e, 'h1099a, 'h1086e, 'h1087e, 'h1099b, 'h1088e, 'h1089e, 'h1099c, 'h108ae, 'h103bc, 'h108be, 'h1099d, 'h108ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1099e, 'h10b9e, 'h106ee, 'h106fe, 'h1099f, 'h1070e, 'h1071e, 'h109a0, 'h1072e, 'h1073e, 'h109a1, 'h1074e, 'h1075e, 'h109a2, 'h103bc, 'h1076e, 'h1077e, 'h109a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078e, 'h10b9e, 'h1079e, 'h109a4, 'h107ae, 'h107be, 'h109a5, 'h107ce, 'h107de, 'h109a6, 'h107ee, 'h107fe, 'h109a7, 'h1080e, 'h103bc, 'h1081e, 'h109a8, 'h1082e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083e, 'h109a9, 'h10b9e, 'h1084e, 'h1085e, 'h109aa, 'h1086e, 'h1087e, 'h109ab, 'h1088e, 'h1089e, 'h109ac, 'h108ae, 'h108be, 'h109ad, 'h103bc, 'h108ce, 'h106de, 'h109ae, 'h10bae, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ee, 'h106fe, 'h109af, 'h1070e, 'h1071e, 'h109b0, 'h1072e, 'h1073e, 'h109b1, 'h1074e, 'h1075e, 'h109b2, 'h1076e, 'h103bc, 'h1077e, 'h109b3, 'h1078e, 'h10bae, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079e, 'h109b4, 'h107ae, 'h107be, 'h109b5, 'h107ce, 'h107de, 'h109b6, 'h107ee, 'h107fe, 'h109b7, 'h1080e, 'h1081e, 'h109b8, 'h103bc, 'h1082e, 'h1083e, 'h109b9, 'h10bae, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084e, 'h1085e, 'h109ba, 'h1086e, 'h1087e, 'h109bb, 'h1088e, 'h1089e, 'h109bc, 'h108ae, 'h108be, 'h109bd, 'h108ce, 'h103bc, 'h106de, 'h109be, 'h10bbe, 'h106ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fe, 'h109bf, 'h1070e, 'h1071e, 'h109c0, 'h1072e, 'h1073e, 'h109c1, 'h1074e, 'h1075e, 'h109c2, 'h1076e, 'h1077e, 'h109c3, 'h103bc, 'h1078e, 'h10bbe, 'h1079e, 'h109c4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ae, 'h107be, 'h109c5, 'h107ce, 'h107de, 'h109c6, 'h107ee, 'h107fe, 'h109c7, 'h1080e, 'h1081e, 'h109c8, 'h1082e, 'h103bc, 'h1083e, 'h109c9, 'h10bbe, 'h1084e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085e, 'h109ca, 'h1086e, 'h1087e, 'h109cb, 'h1088e, 'h1089e, 'h109cc, 'h108ae, 'h108be, 'h109cd, 'h108ce, 'h106de, 'h109ce, 'h10bce, 'h103bc, 'h106ee, 'h106fe, 'h109cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070e, 'h1071e, 'h109d0, 'h1072e, 'h1073e, 'h109d1, 'h1074e, 'h1075e, 'h109d2, 'h1076e, 'h1077e, 'h109d3, 'h1078e, 'h10bce, 'h103bc, 'h1079e, 'h109d4, 'h107ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h107be, 'h109d5, 'h107ce, 'h107de, 'h109d6, 'h107ee, 'h107fe, 'h109d7, 'h1080e, 'h1081e, 'h109d8, 'h1082e, 'h1083e, 'h109d9, 'h10bce, 'h103bc, 'h1084e, 'h1085e, 'h109da, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086e, 'h1087e, 'h109db, 'h1088e, 'h1089e, 'h109dc, 'h108ae, 'h108be, 'h109dd, 'h108ce, 'h106de, 'h109de, 'h10bde, 'h106ee, 'h103bc, 'h106fe, 'h109df, 'h1070e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071e, 'h109e0, 'h1072e, 'h1073e, 'h109e1, 'h1074e, 'h1075e, 'h109e2, 'h1076e, 'h1077e, 'h109e3, 'h1078e, 'h10bde, 'h1079e, 'h109e4, 'h103bc, 'h107ae, 'h107be, 'h109e5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ce, 'h107de, 'h109e6, 'h107ee, 'h107fe, 'h109e7, 'h1080e, 'h1081e, 'h109e8, 'h1082e, 'h1083e, 'h109e9, 'h10bde, 'h1084e, 'h103bc, 'h1085e, 'h109ea, 'h1086e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087e, 'h109eb, 'h1088e, 'h1089e, 'h109ec, 'h108ae, 'h108be, 'h109ed, 'h108ce, 'h106de, 'h109ee, 'h10bee, 'h106ee, 'h106fe, 'h109ef, 'h103bc, 'h1070e, 'h1071e, 'h109f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072e, 'h1073e, 'h109f1, 'h1074e, 'h1075e, 'h109f2, 'h1076e, 'h1077e, 'h109f3, 'h1078e, 'h10bee, 'h1079e, 'h109f4, 'h107ae, 'h103bc, 'h107be, 'h109f5, 'h107ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h107de, 'h109f6, 'h107ee, 'h107fe, 'h109f7, 'h1080e, 'h1081e, 'h109f8, 'h1082e, 'h1083e, 'h109f9, 'h10bee, 'h1084e, 'h1085e, 'h109fa, 'h103bc, 'h1086e, 'h1087e, 'h109fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088e, 'h1089e, 'h109fc, 'h108ae, 'h108be, 'h109fd, 'h108ce, 'h106de, 'h109fe, 'h10bfe, 'h106ee, 'h106fe, 'h109ff, 'h1070e, 'h103bc, 'h1071e, 'h10a00, 'h1072e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073e, 'h10a01, 'h1074e, 'h1075e, 'h10a02, 'h1076e, 'h1077e, 'h10a03, 'h1078e, 'h10bfe, 'h1079e, 'h10a04, 'h107ae, 'h107be, 'h10a05, 'h103bc, 'h107ce, 'h107de, 'h10a06, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ee, 'h107fe, 'h10a07, 'h1080e, 'h1081e, 'h10a08, 'h1082e, 'h1083e, 'h10a09, 'h10bfe, 'h1084e, 'h1085e, 'h10a0a, 'h1086e, 'h103bc, 'h1087e, 'h10a0b, 'h1088e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089e, 'h10a0c, 'h108ae, 'h108be, 'h10a0d, 'h108ce, 'h106de, 'h10a0e, 'h10c0e, 'h106ee, 'h106fe, 'h10a0f, 'h1070e, 'h1071e, 'h10a10, 'h103bc, 'h1072e, 'h1073e, 'h10a11, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074e, 'h1075e, 'h10a12, 'h1076e, 'h1077e, 'h10a13, 'h1078e, 'h10c0e, 'h1079e, 'h10a14, 'h107ae, 'h107be, 'h10a15, 'h107ce, 'h103bc, 'h107de, 'h10a16, 'h107ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fe, 'h10a17, 'h1080e, 'h1081e, 'h10a18, 'h1082e, 'h1083e, 'h10a19, 'h10c0e, 'h1084e, 'h1085e, 'h10a1a, 'h1086e, 'h1087e, 'h10a1b, 'h103bc, 'h1088e, 'h1089e, 'h10a1c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ae, 'h108be, 'h10a1d, 'h108ce, 'h106de, 'h10a1e, 'h10c1e, 'h106ee, 'h106fe, 'h10a1f, 'h1070e, 'h1071e, 'h10a20, 'h1072e, 'h103bc, 'h1073e, 'h10a21, 'h1074e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075e, 'h10a22, 'h1076e, 'h1077e, 'h10a23, 'h1078e, 'h10c1e, 'h1079e, 'h10a24, 'h107ae, 'h107be, 'h10a25, 'h107ce, 'h107de, 'h10a26, 'h103bc, 'h107ee, 'h107fe, 'h10a27, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080e, 'h1081e, 'h10a28, 'h1082e, 'h1083e, 'h10a29, 'h10c1e, 'h1084e, 'h1085e, 'h10a2a, 'h1086e, 'h1087e, 'h10a2b, 'h1088e, 'h103bc, 'h1089e, 'h10a2c, 'h108ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h108be, 'h10a2d, 'h108ce, 'h106de, 'h10a2e, 'h10c2e, 'h106ee, 'h106fe, 'h10a2f, 'h1070e, 'h1071e, 'h10a30, 'h1072e, 'h1073e, 'h10a31, 'h103bc, 'h1074e, 'h1075e, 'h10a32, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076e, 'h1077e, 'h10a33, 'h1078e, 'h10c2e, 'h1079e, 'h10a34, 'h107ae, 'h107be, 'h10a35, 'h107ce, 'h107de, 'h10a36, 'h107ee, 'h103bc, 'h107fe, 'h10a37, 'h1080e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081e, 'h10a38, 'h1082e, 'h1083e, 'h10a39, 'h10c2e, 'h1084e, 'h1085e, 'h10a3a, 'h1086e, 'h1087e, 'h10a3b, 'h1088e, 'h1089e, 'h10a3c, 'h103bc, 'h108ae, 'h108be, 'h10a3d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ce, 'h106de, 'h10a3e, 'h10c3e, 'h106ee, 'h106fe, 'h10a3f, 'h1070e, 'h1071e, 'h10a40, 'h1072e, 'h1073e, 'h10a41, 'h1074e, 'h103bc, 'h1075e, 'h10a42, 'h1076e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077e, 'h10a43, 'h1078e, 'h10c3e, 'h1079e, 'h10a44, 'h107ae, 'h107be, 'h10a45, 'h107ce, 'h107de, 'h10a46, 'h107ee, 'h107fe, 'h10a47, 'h103bc, 'h1080e, 'h1081e, 'h10a48, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082e, 'h1083e, 'h10a49, 'h10c3e, 'h1084e, 'h1085e, 'h10a4a, 'h1086e, 'h1087e, 'h10a4b, 'h1088e, 'h1089e, 'h10a4c, 'h108ae, 'h103bc, 'h108be, 'h10a4d, 'h108ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h10a4e, 'h10c4e, 'h106ee, 'h106fe, 'h10a4f, 'h1070e, 'h1071e, 'h10a50, 'h1072e, 'h1073e, 'h10a51, 'h1074e, 'h1075e, 'h10a52, 'h103bc, 'h1076e, 'h1077e, 'h10a53, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078e, 'h10c4e, 'h1079e, 'h10a54, 'h107ae, 'h107be, 'h10a55, 'h107ce, 'h107de, 'h10a56, 'h107ee, 'h107fe, 'h10a57, 'h1080e, 'h103bc, 'h1081e, 'h10a58, 'h1082e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083e, 'h10a59, 'h10c4e, 'h1084e, 'h1085e, 'h10a5a, 'h1086e, 'h1087e, 'h10a5b, 'h1088e, 'h1089e, 'h10a5c, 'h108ae, 'h108be, 'h10a5d, 'h103bc, 'h108ce, 'h106de, 'h10a5e, 'h10c5e, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ee, 'h106fe, 'h10a5f, 'h1070e, 'h1071e, 'h10a60, 'h1072e, 'h1073e, 'h10a61, 'h1074e, 'h1075e, 'h10a62, 'h1076e, 'h103bc, 'h1077e, 'h10a63, 'h1078e, 'h10c5e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079e, 'h10a64, 'h107ae, 'h107be, 'h10a65, 'h107ce, 'h107de, 'h10a66, 'h107ee, 'h107fe, 'h10a67, 'h1080e, 'h1081e, 'h10a68, 'h103bc, 'h1082e, 'h1083e, 'h10a69, 'h10c5e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084e, 'h1085e, 'h10a6a, 'h1086e, 'h1087e, 'h10a6b, 'h1088e, 'h1089e, 'h10a6c, 'h108ae, 'h108be, 'h10a6d, 'h108ce, 'h103bc, 'h106de, 'h10a6e, 'h10c6e, 'h106ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h106fe, 'h10a6f, 'h1070e, 'h1071e, 'h10a70, 'h1072e, 'h1073e, 'h10a71, 'h1074e, 'h1075e, 'h10a72, 'h1076e, 'h1077e, 'h10a73, 'h103bc, 'h1078e, 'h10c6e, 'h1079e, 'h10a74, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ae, 'h107be, 'h10a75, 'h107ce, 'h107de, 'h10a76, 'h107ee, 'h107fe, 'h10a77, 'h1080e, 'h1081e, 'h10a78, 'h1082e, 'h103bc, 'h1083e, 'h10a79, 'h10c6e, 'h1084e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085e, 'h10a7a, 'h1086e, 'h1087e, 'h10a7b, 'h1088e, 'h1089e, 'h10a7c, 'h108ae, 'h108be, 'h10a7d, 'h108ce, 'h106de, 'h10a7e, 'h10c7e, 'h103bc, 'h106ee, 'h106fe, 'h10a7f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070e, 'h1071e, 'h10a80, 'h1072e, 'h1073e, 'h10a81, 'h1074e, 'h1075e, 'h10a82, 'h1076e, 'h1077e, 'h10a83, 'h1078e, 'h10c7e, 'h103bc, 'h1079e, 'h10a84, 'h107ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h107be, 'h10a85, 'h107ce, 'h107de, 'h10a86, 'h107ee, 'h107fe, 'h10a87, 'h1080e, 'h1081e, 'h10a88, 'h1082e, 'h1083e, 'h10a89, 'h10c7e, 'h103bc, 'h1084e, 'h1085e, 'h10a8a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086e, 'h1087e, 'h10a8b, 'h1088e, 'h1089e, 'h10a8c, 'h108ae, 'h108be, 'h10a8d, 'h108ce, 'h106de, 'h10a8e, 'h10c8e, 'h106ee, 'h103bc, 'h106fe, 'h10a8f, 'h1070e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071e, 'h10a90, 'h1072e, 'h1073e, 'h10a91, 'h1074e, 'h1075e, 'h10a92, 'h1076e, 'h1077e, 'h10a93, 'h1078e, 'h10c8e, 'h1079e, 'h10a94, 'h103bc, 'h107ae, 'h107be, 'h10a95, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ce, 'h107de, 'h10a96, 'h107ee, 'h107fe, 'h10a97, 'h1080e, 'h1081e, 'h10a98, 'h1082e, 'h1083e, 'h10a99, 'h10c8e, 'h1084e, 'h103bc, 'h1085e, 'h10a9a, 'h1086e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087e, 'h10a9b, 'h1088e, 'h1089e, 'h10a9c, 'h108ae, 'h108be, 'h10a9d, 'h108ce, 'h106de, 'h10a9e, 'h10c9e, 'h106ee, 'h106fe, 'h10a9f, 'h103bc, 'h1070e, 'h1071e, 'h10aa0, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072e, 'h1073e, 'h10aa1, 'h1074e, 'h1075e, 'h10aa2, 'h1076e, 'h1077e, 'h10aa3, 'h1078e, 'h10c9e, 'h1079e, 'h10aa4, 'h107ae, 'h103bc, 'h107be, 'h10aa5, 'h107ce, 'h21f8e, 'h21f8f, 'h21f8d, 'h107de, 'h10aa6, 'h107ee, 'h107fe, 'h10aa7, 'h1080e, 'h1081e, 'h10aa8, 'h1082e, 'h1083e, 'h10aa9, 'h10c9e, 'h1084e, 'h1085e, 'h10aaa, 'h103bc, 'h1086e, 'h1087e, 'h10aab, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088e, 'h1089e, 'h10aac, 'h108ae, 'h108be, 'h10aad, 'h108ce, 'h106de, 'h10aae, 'h10cae, 'h106ee, 'h106fe, 'h10aaf, 'h1070e, 'h103bc, 'h1071e, 'h10ab0, 'h1072e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073e, 'h10ab1, 'h1074e, 'h1075e, 'h10ab2, 'h1076e, 'h1077e, 'h10ab3, 'h1078e, 'h10cae, 'h1079e, 'h10ab4, 'h107ae, 'h107be, 'h10ab5, 'h103bc, 'h107ce, 'h107de, 'h10ab6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ee, 'h107fe, 'h10ab7, 'h1080e, 'h1081e, 'h10ab8, 'h1082e, 'h1083e, 'h10ab9, 'h10cae, 'h1084e, 'h1085e, 'h10aba, 'h1086e, 'h103bc, 'h1087e, 'h10abb, 'h1088e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089e, 'h10abc, 'h108ae, 'h108be, 'h10abd, 'h108ce, 'h106de, 'h10abe, 'h10cbe, 'h106ee, 'h106fe, 'h10abf, 'h1070e, 'h1071e, 'h10ac0, 'h103bc, 'h1072e, 'h1073e, 'h10ac1, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074e, 'h1075e, 'h10ac2, 'h1076e, 'h1077e, 'h10ac3, 'h1078e, 'h10cbe, 'h1079e, 'h10ac4, 'h107ae, 'h107be, 'h10ac5, 'h107ce, 'h103bc, 'h107de, 'h10ac6, 'h107ee, 'h21f8e, 'h21f8f, 'h21f8d, 'h107fe, 'h10ac7, 'h1080e, 'h1081e, 'h10ac8, 'h1082e, 'h1083e, 'h10ac9, 'h10cbe, 'h1084e, 'h1085e, 'h10aca, 'h1086e, 'h1087e, 'h10acb, 'h103bc, 'h1088e, 'h1089e, 'h10acc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108ae, 'h108be, 'h10acd, 'h108ce, 'h106de, 'h10ace, 'h10cce, 'h106ee, 'h106fe, 'h10acf, 'h1070e, 'h1071e, 'h10ad0, 'h1072e, 'h103bc, 'h1073e, 'h10ad1, 'h1074e, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075e, 'h10ad2, 'h1076e, 'h1077e, 'h10ad3, 'h1078e, 'h10cce, 'h1079e, 'h10ad4, 'h107ae, 'h107be, 'h10ad5, 'h107ce, 'h107de, 'h10ad6, 'h103bc, 'h107ee, 'h107fe, 'h10ad7, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080e, 'h1081e, 'h10ad8, 'h1082e, 'h1083e, 'h10ad9, 'h10cce, 'h1084e, 'h1085e, 'h10ada, 'h1086e, 'h1087e, 'h10adb, 'h1088e, 'h103bc, 'h1089e, 'h10adc, 'h108ae, 'h21f8e, 'h21f8f, 'h21f8d, 'h108be, 'h10add, 'h108ce, 'h106df, 'h108de, 'h10adf, 'h106ef, 'h106ff, 'h108df, 'h1070f, 'h1071f, 'h108e0, 'h1072f, 'h1073f, 'h108e1, 'h103bc, 'h1074f, 'h1075f, 'h108e2, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076f, 'h1077f, 'h108e3, 'h1078f, 'h10adf, 'h1079f, 'h108e4, 'h107af, 'h107bf, 'h108e5, 'h107cf, 'h107df, 'h108e6, 'h107ef, 'h103bc, 'h107ff, 'h108e7, 'h1080f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081f, 'h108e8, 'h1082f, 'h1083f, 'h108e9, 'h10adf, 'h1084f, 'h1085f, 'h108ea, 'h1086f, 'h1087f, 'h108eb, 'h1088f, 'h1089f, 'h108ec, 'h103bc, 'h108af, 'h108bf, 'h108ed, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cf, 'h106df, 'h108ee, 'h10aef, 'h106ef, 'h106ff, 'h108ef, 'h1070f, 'h1071f, 'h108f0, 'h1072f, 'h1073f, 'h108f1, 'h1074f, 'h103bc, 'h1075f, 'h108f2, 'h1076f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077f, 'h108f3, 'h1078f, 'h10aef, 'h1079f, 'h108f4, 'h107af, 'h107bf, 'h108f5, 'h107cf, 'h107df, 'h108f6, 'h107ef, 'h107ff, 'h108f7, 'h103bc, 'h1080f, 'h1081f, 'h108f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082f, 'h1083f, 'h108f9, 'h10aef, 'h1084f, 'h1085f, 'h108fa, 'h1086f, 'h1087f, 'h108fb, 'h1088f, 'h1089f, 'h108fc, 'h108af, 'h103bc, 'h108bf, 'h108fd, 'h108cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h108fe, 'h10aff, 'h106ef, 'h106ff, 'h108ff, 'h1070f, 'h1071f, 'h10900, 'h1072f, 'h1073f, 'h10901, 'h1074f, 'h1075f, 'h10902, 'h103bc, 'h1076f, 'h1077f, 'h10903, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078f, 'h10aff, 'h1079f, 'h10904, 'h107af, 'h107bf, 'h10905, 'h107cf, 'h107df, 'h10906, 'h107ef, 'h107ff, 'h10907, 'h1080f, 'h103bc, 'h1081f, 'h10908, 'h1082f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083f, 'h10909, 'h10aff, 'h1084f, 'h1085f, 'h1090a, 'h1086f, 'h1087f, 'h1090b, 'h1088f, 'h1089f, 'h1090c, 'h108af, 'h108bf, 'h1090d, 'h103bc, 'h108cf, 'h106df, 'h1090e, 'h10b0f, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ef, 'h106ff, 'h1090f, 'h1070f, 'h1071f, 'h10910, 'h1072f, 'h1073f, 'h10911, 'h1074f, 'h1075f, 'h10912, 'h1076f, 'h103bc, 'h1077f, 'h10913, 'h1078f, 'h10b0f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079f, 'h10914, 'h107af, 'h107bf, 'h10915, 'h107cf, 'h107df, 'h10916, 'h107ef, 'h107ff, 'h10917, 'h1080f, 'h1081f, 'h10918, 'h103bc, 'h1082f, 'h1083f, 'h10919, 'h10b0f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084f, 'h1085f, 'h1091a, 'h1086f, 'h1087f, 'h1091b, 'h1088f, 'h1089f, 'h1091c, 'h108af, 'h108bf, 'h1091d, 'h108cf, 'h103bc, 'h106df, 'h1091e, 'h10b1f, 'h106ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ff, 'h1091f, 'h1070f, 'h1071f, 'h10920, 'h1072f, 'h1073f, 'h10921, 'h1074f, 'h1075f, 'h10922, 'h1076f, 'h1077f, 'h10923, 'h103bc, 'h1078f, 'h10b1f, 'h1079f, 'h10924, 'h21f8e, 'h21f8f, 'h21f8d, 'h107af, 'h107bf, 'h10925, 'h107cf, 'h107df, 'h10926, 'h107ef, 'h107ff, 'h10927, 'h1080f, 'h1081f, 'h10928, 'h1082f, 'h103bc, 'h1083f, 'h10929, 'h10b1f, 'h1084f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085f, 'h1092a, 'h1086f, 'h1087f, 'h1092b, 'h1088f, 'h1089f, 'h1092c, 'h108af, 'h108bf, 'h1092d, 'h108cf, 'h106df, 'h1092e, 'h10b2f, 'h103bc, 'h106ef, 'h106ff, 'h1092f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070f, 'h1071f, 'h10930, 'h1072f, 'h1073f, 'h10931, 'h1074f, 'h1075f, 'h10932, 'h1076f, 'h1077f, 'h10933, 'h1078f, 'h10b2f, 'h103bc, 'h1079f, 'h10934, 'h107af, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bf, 'h10935, 'h107cf, 'h107df, 'h10936, 'h107ef, 'h107ff, 'h10937, 'h1080f, 'h1081f, 'h10938, 'h1082f, 'h1083f, 'h10939, 'h10b2f, 'h103bc, 'h1084f, 'h1085f, 'h1093a, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086f, 'h1087f, 'h1093b, 'h1088f, 'h1089f, 'h1093c, 'h108af, 'h108bf, 'h1093d, 'h108cf, 'h106df, 'h1093e, 'h10b3f, 'h106ef, 'h103bc, 'h106ff, 'h1093f, 'h1070f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071f, 'h10940, 'h1072f, 'h1073f, 'h10941, 'h1074f, 'h1075f, 'h10942, 'h1076f, 'h1077f, 'h10943, 'h1078f, 'h10b3f, 'h1079f, 'h10944, 'h103bc, 'h107af, 'h107bf, 'h10945, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cf, 'h107df, 'h10946, 'h107ef, 'h107ff, 'h10947, 'h1080f, 'h1081f, 'h10948, 'h1082f, 'h1083f, 'h10949, 'h10b3f, 'h1084f, 'h103bc, 'h1085f, 'h1094a, 'h1086f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087f, 'h1094b, 'h1088f, 'h1089f, 'h1094c, 'h108af, 'h108bf, 'h1094d, 'h108cf, 'h106df, 'h1094e, 'h10b4f, 'h106ef, 'h106ff, 'h1094f, 'h103bc, 'h1070f, 'h1071f, 'h10950, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072f, 'h1073f, 'h10951, 'h1074f, 'h1075f, 'h10952, 'h1076f, 'h1077f, 'h10953, 'h1078f, 'h10b4f, 'h1079f, 'h10954, 'h107af, 'h103bc, 'h107bf, 'h10955, 'h107cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h107df, 'h10956, 'h107ef, 'h107ff, 'h10957, 'h1080f, 'h1081f, 'h10958, 'h1082f, 'h1083f, 'h10959, 'h10b4f, 'h1084f, 'h1085f, 'h1095a, 'h103bc, 'h1086f, 'h1087f, 'h1095b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088f, 'h1089f, 'h1095c, 'h108af, 'h108bf, 'h1095d, 'h108cf, 'h106df, 'h1095e, 'h10b5f, 'h106ef, 'h106ff, 'h1095f, 'h1070f, 'h103bc, 'h1071f, 'h10960, 'h1072f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073f, 'h10961, 'h1074f, 'h1075f, 'h10962, 'h1076f, 'h1077f, 'h10963, 'h1078f, 'h10b5f, 'h1079f, 'h10964, 'h107af, 'h107bf, 'h10965, 'h103bc, 'h107cf, 'h107df, 'h10966, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ef, 'h107ff, 'h10967, 'h1080f, 'h1081f, 'h10968, 'h1082f, 'h1083f, 'h10969, 'h10b5f, 'h1084f, 'h1085f, 'h1096a, 'h1086f, 'h103bc, 'h1087f, 'h1096b, 'h1088f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089f, 'h1096c, 'h108af, 'h108bf, 'h1096d, 'h108cf, 'h106df, 'h1096e, 'h10b6f, 'h106ef, 'h106ff, 'h1096f, 'h1070f, 'h1071f, 'h10970, 'h103bc, 'h1072f, 'h1073f, 'h10971, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074f, 'h1075f, 'h10972, 'h1076f, 'h1077f, 'h10973, 'h1078f, 'h10b6f, 'h1079f, 'h10974, 'h107af, 'h107bf, 'h10975, 'h107cf, 'h103bc, 'h107df, 'h10976, 'h107ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ff, 'h10977, 'h1080f, 'h1081f, 'h10978, 'h1082f, 'h1083f, 'h10979, 'h10b6f, 'h1084f, 'h1085f, 'h1097a, 'h1086f, 'h1087f, 'h1097b, 'h103bc, 'h1088f, 'h1089f, 'h1097c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108af, 'h108bf, 'h1097d, 'h108cf, 'h106df, 'h1097e, 'h10b7f, 'h106ef, 'h106ff, 'h1097f, 'h1070f, 'h1071f, 'h10980, 'h1072f, 'h103bc, 'h1073f, 'h10981, 'h1074f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075f, 'h10982, 'h1076f, 'h1077f, 'h10983, 'h1078f, 'h10b7f, 'h1079f, 'h10984, 'h107af, 'h107bf, 'h10985, 'h107cf, 'h107df, 'h10986, 'h103bc, 'h107ef, 'h107ff, 'h10987, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080f, 'h1081f, 'h10988, 'h1082f, 'h1083f, 'h10989, 'h10b7f, 'h1084f, 'h1085f, 'h1098a, 'h1086f, 'h1087f, 'h1098b, 'h1088f, 'h103bc, 'h1089f, 'h1098c, 'h108af, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bf, 'h1098d, 'h108cf, 'h106df, 'h1098e, 'h10b8f, 'h106ef, 'h106ff, 'h1098f, 'h1070f, 'h1071f, 'h10990, 'h1072f, 'h1073f, 'h10991, 'h103bc, 'h1074f, 'h1075f, 'h10992, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076f, 'h1077f, 'h10993, 'h1078f, 'h10b8f, 'h1079f, 'h10994, 'h107af, 'h107bf, 'h10995, 'h107cf, 'h107df, 'h10996, 'h107ef, 'h103bc, 'h107ff, 'h10997, 'h1080f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081f, 'h10998, 'h1082f, 'h1083f, 'h10999, 'h10b8f, 'h1084f, 'h1085f, 'h1099a, 'h1086f, 'h1087f, 'h1099b, 'h1088f, 'h1089f, 'h1099c, 'h103bc, 'h108af, 'h108bf, 'h1099d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cf, 'h106df, 'h1099e, 'h10b9f, 'h106ef, 'h106ff, 'h1099f, 'h1070f, 'h1071f, 'h109a0, 'h1072f, 'h1073f, 'h109a1, 'h1074f, 'h103bc, 'h1075f, 'h109a2, 'h1076f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077f, 'h109a3, 'h1078f, 'h10b9f, 'h1079f, 'h109a4, 'h107af, 'h107bf, 'h109a5, 'h107cf, 'h107df, 'h109a6, 'h107ef, 'h107ff, 'h109a7, 'h103bc, 'h1080f, 'h1081f, 'h109a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082f, 'h1083f, 'h109a9, 'h10b9f, 'h1084f, 'h1085f, 'h109aa, 'h1086f, 'h1087f, 'h109ab, 'h1088f, 'h1089f, 'h109ac, 'h108af, 'h103bc, 'h108bf, 'h109ad, 'h108cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h109ae, 'h10baf, 'h106ef, 'h106ff, 'h109af, 'h1070f, 'h1071f, 'h109b0, 'h1072f, 'h1073f, 'h109b1, 'h1074f, 'h1075f, 'h109b2, 'h103bc, 'h1076f, 'h1077f, 'h109b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1078f, 'h10baf, 'h1079f, 'h109b4, 'h107af, 'h107bf, 'h109b5, 'h107cf, 'h107df, 'h109b6, 'h107ef, 'h107ff, 'h109b7, 'h1080f, 'h103bc, 'h1081f, 'h109b8, 'h1082f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1083f, 'h109b9, 'h10baf, 'h1084f, 'h1085f, 'h109ba, 'h1086f, 'h1087f, 'h109bb, 'h1088f, 'h1089f, 'h109bc, 'h108af, 'h108bf, 'h109bd, 'h103bc, 'h108cf, 'h106df, 'h109be, 'h10bbf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ef, 'h106ff, 'h109bf, 'h1070f, 'h1071f, 'h109c0, 'h1072f, 'h1073f, 'h109c1, 'h1074f, 'h1075f, 'h109c2, 'h1076f, 'h103bc, 'h1077f, 'h109c3, 'h1078f, 'h10bbf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1079f, 'h109c4, 'h107af, 'h107bf, 'h109c5, 'h107cf, 'h107df, 'h109c6, 'h107ef, 'h107ff, 'h109c7, 'h1080f, 'h1081f, 'h109c8, 'h103bc, 'h1082f, 'h1083f, 'h109c9, 'h10bbf, 'h21f8e, 'h21f8f, 'h21f8d, 'h1084f, 'h1085f, 'h109ca, 'h1086f, 'h1087f, 'h109cb, 'h1088f, 'h1089f, 'h109cc, 'h108af, 'h108bf, 'h109cd, 'h108cf, 'h103bc, 'h106df, 'h109ce, 'h10bcf, 'h106ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h106ff, 'h109cf, 'h1070f, 'h1071f, 'h109d0, 'h1072f, 'h1073f, 'h109d1, 'h1074f, 'h1075f, 'h109d2, 'h1076f, 'h1077f, 'h109d3, 'h103bc, 'h1078f, 'h10bcf, 'h1079f, 'h109d4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107af, 'h107bf, 'h109d5, 'h107cf, 'h107df, 'h109d6, 'h107ef, 'h107ff, 'h109d7, 'h1080f, 'h1081f, 'h109d8, 'h1082f, 'h103bc, 'h1083f, 'h109d9, 'h10bcf, 'h1084f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1085f, 'h109da, 'h1086f, 'h1087f, 'h109db, 'h1088f, 'h1089f, 'h109dc, 'h108af, 'h108bf, 'h109dd, 'h108cf, 'h106df, 'h109de, 'h10bdf, 'h103bc, 'h106ef, 'h106ff, 'h109df, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070f, 'h1071f, 'h109e0, 'h1072f, 'h1073f, 'h109e1, 'h1074f, 'h1075f, 'h109e2, 'h1076f, 'h1077f, 'h109e3, 'h1078f, 'h10bdf, 'h103bc, 'h1079f, 'h109e4, 'h107af, 'h21f8e, 'h21f8f, 'h21f8d, 'h107bf, 'h109e5, 'h107cf, 'h107df, 'h109e6, 'h107ef, 'h107ff, 'h109e7, 'h1080f, 'h1081f, 'h109e8, 'h1082f, 'h1083f, 'h109e9, 'h10bdf, 'h103bc, 'h1084f, 'h1085f, 'h109ea, 'h21f8e, 'h21f8f, 'h21f8d, 'h1086f, 'h1087f, 'h109eb, 'h1088f, 'h1089f, 'h109ec, 'h108af, 'h108bf, 'h109ed, 'h108cf, 'h106df, 'h109ee, 'h10bef, 'h106ef, 'h103bc, 'h106ff, 'h109ef, 'h1070f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1071f, 'h109f0, 'h1072f, 'h1073f, 'h109f1, 'h1074f, 'h1075f, 'h109f2, 'h1076f, 'h1077f, 'h109f3, 'h1078f, 'h10bef, 'h1079f, 'h109f4, 'h103bc, 'h107af, 'h107bf, 'h109f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107cf, 'h107df, 'h109f6, 'h107ef, 'h107ff, 'h109f7, 'h1080f, 'h1081f, 'h109f8, 'h1082f, 'h1083f, 'h109f9, 'h10bef, 'h1084f, 'h103bc, 'h1085f, 'h109fa, 'h1086f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1087f, 'h109fb, 'h1088f, 'h1089f, 'h109fc, 'h108af, 'h108bf, 'h109fd, 'h108cf, 'h106df, 'h109fe, 'h10bff, 'h106ef, 'h106ff, 'h109ff, 'h103bc, 'h1070f, 'h1071f, 'h10a00, 'h21f8e, 'h21f8f, 'h21f8d, 'h1072f, 'h1073f, 'h10a01, 'h1074f, 'h1075f, 'h10a02, 'h1076f, 'h1077f, 'h10a03, 'h1078f, 'h10bff, 'h1079f, 'h10a04, 'h107af, 'h103bc, 'h107bf, 'h10a05, 'h107cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h107df, 'h10a06, 'h107ef, 'h107ff, 'h10a07, 'h1080f, 'h1081f, 'h10a08, 'h1082f, 'h1083f, 'h10a09, 'h10bff, 'h1084f, 'h1085f, 'h10a0a, 'h103bc, 'h1086f, 'h1087f, 'h10a0b, 'h21f8e, 'h21f8f, 'h21f8d, 'h1088f, 'h1089f, 'h10a0c, 'h108af, 'h108bf, 'h10a0d, 'h108cf, 'h106df, 'h10a0e, 'h10c0f, 'h106ef, 'h106ff, 'h10a0f, 'h1070f, 'h103bc, 'h1071f, 'h10a10, 'h1072f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073f, 'h10a11, 'h1074f, 'h1075f, 'h10a12, 'h1076f, 'h1077f, 'h10a13, 'h1078f, 'h10c0f, 'h1079f, 'h10a14, 'h107af, 'h107bf, 'h10a15, 'h103bc, 'h107cf, 'h107df, 'h10a16, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ef, 'h107ff, 'h10a17, 'h1080f, 'h1081f, 'h10a18, 'h1082f, 'h1083f, 'h10a19, 'h10c0f, 'h1084f, 'h1085f, 'h10a1a, 'h1086f, 'h103bc, 'h1087f, 'h10a1b, 'h1088f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1089f, 'h10a1c, 'h108af, 'h108bf, 'h10a1d, 'h108cf, 'h106df, 'h10a1e, 'h10c1f, 'h106ef, 'h106ff, 'h10a1f, 'h1070f, 'h1071f, 'h10a20, 'h103bc, 'h1072f, 'h1073f, 'h10a21, 'h21f8e, 'h21f8f, 'h21f8d, 'h1074f, 'h1075f, 'h10a22, 'h1076f, 'h1077f, 'h10a23, 'h1078f, 'h10c1f, 'h1079f, 'h10a24, 'h107af, 'h107bf, 'h10a25, 'h107cf, 'h103bc, 'h107df, 'h10a26, 'h107ef, 'h21f8e, 'h21f8f, 'h21f8d, 'h107ff, 'h10a27, 'h1080f, 'h1081f, 'h10a28, 'h1082f, 'h1083f, 'h10a29, 'h10c1f, 'h1084f, 'h1085f, 'h10a2a, 'h1086f, 'h1087f, 'h10a2b, 'h103bc, 'h1088f, 'h1089f, 'h10a2c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108af, 'h108bf, 'h10a2d, 'h108cf, 'h106df, 'h10a2e, 'h10c2f, 'h106ef, 'h106ff, 'h10a2f, 'h1070f, 'h1071f, 'h10a30, 'h1072f, 'h103bc, 'h1073f, 'h10a31, 'h1074f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1075f, 'h10a32, 'h1076f, 'h1077f, 'h10a33, 'h1078f, 'h10c2f, 'h1079f, 'h10a34, 'h107af, 'h107bf, 'h10a35, 'h107cf, 'h107df, 'h10a36, 'h103bc, 'h107ef, 'h107ff, 'h10a37, 'h21f8e, 'h21f8f, 'h21f8d, 'h1080f, 'h1081f, 'h10a38, 'h1082f, 'h1083f, 'h10a39, 'h10c2f, 'h1084f, 'h1085f, 'h10a3a, 'h1086f, 'h1087f, 'h10a3b, 'h1088f, 'h103bc, 'h1089f, 'h10a3c, 'h108af, 'h21f8e, 'h21f8f, 'h21f8d, 'h108bf, 'h10a3d, 'h108cf, 'h106df, 'h10a3e, 'h10c3f, 'h106ef, 'h106ff, 'h10a3f, 'h1070f, 'h1071f, 'h10a40, 'h1072f, 'h1073f, 'h10a41, 'h103bc, 'h1074f, 'h1075f, 'h10a42, 'h21f8e, 'h21f8f, 'h21f8d, 'h1076f, 'h1077f, 'h10a43, 'h1078f, 'h10c3f, 'h1079f, 'h10a44, 'h107af, 'h107bf, 'h10a45, 'h107cf, 'h107df, 'h10a46, 'h107ef, 'h103bc, 'h107ff, 'h10a47, 'h1080f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1081f, 'h10a48, 'h1082f, 'h1083f, 'h10a49, 'h10c3f, 'h1084f, 'h1085f, 'h10a4a, 'h1086f, 'h1087f, 'h10a4b, 'h1088f, 'h1089f, 'h10a4c, 'h103bc, 'h108af, 'h108bf, 'h10a4d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108cf, 'h106df, 'h10a4e, 'h10c4f, 'h106ef, 'h106ff, 'h10a4f, 'h1070f, 'h1071f, 'h10a50, 'h1072f, 'h1073f, 'h10a51, 'h1074f, 'h103bc, 'h1075f, 'h10a52, 'h1076f, 'h21f8e, 'h21f8f, 'h21f8d, 'h1077f, 'h10a53, 'h1078f, 'h10c4f, 'h1079f, 'h10a54, 'h107af, 'h107bf, 'h10a55, 'h107cf, 'h107df, 'h10a56, 'h107ef, 'h107ff, 'h10a57, 'h103bc, 'h1080f, 'h1081f, 'h10a58, 'h21f8e, 'h21f8f, 'h21f8d, 'h1082f, 'h1083f, 'h10a59, 'h10c4f, 'h1084f, 'h1085f, 'h10a5a, 'h1086f, 'h1087f, 'h10a5b, 'h1088f, 'h1089f, 'h10a5c, 'h108af, 'h103bc, 'h108bf, 'h10a5d, 'h108cf, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h10a5e, 'h10c5f, 'h106ef, 'h106ff, 'h10a5f, 'h1070f, 'h1071f, 'h10a60};
	
endpackage
