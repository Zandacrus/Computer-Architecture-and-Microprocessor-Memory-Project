

package LU_PKG_4;
	
	import LU_PKG_3::DATA3;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h100260, 'h100261, 'h100262, 'h100263, 'h1000f0, 'h1000f1, 'h100264, 'h1000f2, 'h10003c, 'h2004f8, 'h100047, 'h100265, 'h1000f3, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000f7, 'h1000f4, 'h10003c, 'h2004f8, 'h100047, 'h1000f5, 'h100172, 'h1000f6, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000f7, 'h10003c, 'h2004f8, 'h100047, 'h100181, 'h1000f4, 'h100182, 'h1000f5, 'h100183, 'h1000f6, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h10003c, 'h2004f8, 'h100047, 'h100190, 'h1000f7, 'h100191, 'h1000f4, 'h100192, 'h1000f5, 'h100193, 'h1000f6, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019d, 'h10003c, 'h2004f8, 'h100047, 'h10019e, 'h10019f, 'h1001a0, 'h1000f7, 'h1001a1, 'h1001a2, 'h1000f4, 'h1000f5, 'h1001a3, 'h1000f6, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h10003c, 'h2004f8, 'h100047, 'h1001af, 'h1001b0, 'h1001b1, 'h1000f7, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1000f4, 'h1000f5, 'h1001b7, 'h1000f6, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h10003c, 'h2004f8, 'h100047, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1000f7, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1000f4, 'h1000f5, 'h1001c7, 'h1000f6, 'h1001c8, 'h1001c9, 'h1001ca, 'h10003c, 'h2004f8, 'h100047, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1000f7, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1000f4, 'h1000f5, 'h1001d7, 'h1000f6, 'h1001d8, 'h10003c, 'h2004f8, 'h100047, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1000f7, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1000f4, 'h1000f5, 'h1001e7, 'h10003c, 'h2004f8, 'h100047, 'h1000f6, 'h1001e8, 'h1001e9, 'h1001ea, 'h1000f7, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1000f4, 'h10003c, 'h2004f8, 'h100047, 'h1001f7, 'h1000f5, 'h1001f8, 'h1000f6, 'h1001f9, 'h1000f7, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h10003c, 'h2004f8, 'h100047, 'h100206, 'h1000f4, 'h100207, 'h1000f5, 'h100208, 'h1000f6, 'h100209, 'h1000f7, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100213, 'h10003c, 'h2004f8, 'h100047, 'h100214, 'h100215, 'h100216, 'h1000f4, 'h100217, 'h1000f5, 'h100218, 'h1000f6, 'h100219, 'h1000f7, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021e, 'h10021f, 'h100220, 'h100221, 'h10003c, 'h2004f8, 'h100047, 'h100222, 'h100223, 'h100224, 'h100225, 'h100227, 'h1000f4, 'h1000f5, 'h100228, 'h1000f6, 'h100229, 'h1000f7, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h10003c, 'h2004f8, 'h100047, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h1000f4, 'h1000f5, 'h100238, 'h1000f6, 'h100239, 'h1000f7, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h10003c, 'h2004f8, 'h100047, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h1000f4, 'h1000f5, 'h100248, 'h1000f6, 'h100249, 'h1000f7, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10003c, 'h2004f8, 'h100047, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h1000f4, 'h1000f5, 'h100258, 'h1000f6, 'h100259, 'h1000f7, 'h10025a, 'h10025b, 'h10025c, 'h10003c, 'h2004f8, 'h100047, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h1000f4, 'h1000f5, 'h100268, 'h1000f6, 'h100269, 'h1000f7, 'h10026a, 'h10003c, 'h2004f8, 'h100047, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000fb, 'h100172, 'h1000f8, 'h1000f9, 'h1000fa, 'h100173, 'h100174, 'h100175, 'h100176, 'h10003c, 'h2004f8, 'h100047, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000fb, 'h100181, 'h100182, 'h1000f8, 'h1000f9, 'h100183, 'h1000fa, 'h100184, 'h10003c, 'h2004f8, 'h100047, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h1000fb, 'h10018f, 'h100190, 'h100191, 'h100193, 'h1000f8, 'h100192, 'h1000f9, 'h10003c, 'h2004f8, 'h100047, 'h1000fa, 'h100194, 'h100195, 'h100197, 'h100196, 'h100198, 'h100199, 'h10019b, 'h10019a, 'h10019c, 'h1000fb, 'h10019d, 'h10019f, 'h10019e, 'h1001a0, 'h1001a2, 'h1001a3, 'h1000f8, 'h10003c, 'h2004f8, 'h100047, 'h1000f9, 'h1000fa, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1000fb, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h10003c, 'h2004f8, 'h100047, 'h1001b6, 'h1001b7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1000fb, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h10003c, 'h2004f8, 'h100047, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1001c8, 'h1001c9, 'h1001ca, 'h1000fb, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h10003c, 'h2004f8, 'h100047, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1001d8, 'h1000fb, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h10003c, 'h2004f8, 'h100047, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1001e8, 'h1000fb, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h10003c, 'h2004f8, 'h100047, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1000f8, 'h1000f9, 'h1000fa, 'h1001f8, 'h1000fb, 'h1001f9, 'h1001fa, 'h1001fb, 'h10003c, 'h2004f8, 'h100047, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100207, 'h1000f8, 'h1000f9, 'h100208, 'h1000fa, 'h100209, 'h1000fb, 'h10003c, 'h2004f8, 'h100047, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100214, 'h100213, 'h100215, 'h100216, 'h100218, 'h1000f8, 'h100217, 'h1000f9, 'h1000fa, 'h10003c, 'h2004f8, 'h100047, 'h100219, 'h1000fb, 'h10021a, 'h10021c, 'h10021b, 'h10021d, 'h10021e, 'h100220, 'h10021f, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h1000f8, 'h1000f9, 'h1000fa, 'h10003c, 'h2004f8, 'h100047, 'h100229, 'h1000fb, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h1000f8, 'h1000f9, 'h1000fa, 'h10003c, 'h2004f8, 'h100047, 'h100239, 'h1000fb, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h1000f8, 'h10003c, 'h2004f8, 'h100047, 'h1000f9, 'h1000fa, 'h100249, 'h1000fb, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h10003c, 'h2004f8, 'h100047, 'h1000f8, 'h1000f9, 'h1000fa, 'h100259, 'h1000fb, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h10003c, 'h2004f8, 'h100047, 'h100267, 'h100268, 'h1000f8, 'h1000f9, 'h1000fa, 'h100269, 'h1000fb, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h1000ff, 'h10003c, 'h2004f8, 'h100047, 'h1000fc, 'h1000fd, 'h100172, 'h1000fe, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h1000ff, 'h10003c, 'h2004f8, 'h100047, 'h100181, 'h1000fc, 'h100182, 'h1000fd, 'h100183, 'h1000fe, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10018e, 'h10018f, 'h10003c, 'h2004f8, 'h100047, 'h100190, 'h1000ff, 'h100191, 'h1000fc, 'h100192, 'h1000fd, 'h100193, 'h1000fe, 'h100194, 'h100195, 'h100196, 'h100197, 'h100198, 'h100199, 'h10019a, 'h10019b, 'h10019c, 'h10019e, 'h10003c, 'h2004f8, 'h100047, 'h10019f, 'h1001a0, 'h1000ff, 'h1001a2, 'h1000fc, 'h1000fd, 'h1001a3, 'h1000fe, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h10003c, 'h2004f8, 'h100047, 'h1001b1, 'h1001b2, 'h1000ff, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1000fc, 'h1000fd, 'h1001b7, 'h1000fe, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h10003c, 'h2004f8, 'h100047, 'h1001bf, 'h1001c0, 'h1000ff, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1000fc, 'h1000fd, 'h1001c7, 'h1000fe, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h10003c, 'h2004f8, 'h100047, 'h1001cd, 'h1001ce, 'h1000ff, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1000fc, 'h1000fd, 'h1001d7, 'h1000fe, 'h1001d8, 'h1001d9, 'h1001da, 'h10003c, 'h2004f8, 'h100047, 'h1001db, 'h1001dc, 'h1000ff, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1000fc, 'h1000fd, 'h1001e7, 'h1000fe, 'h1001e8, 'h10003c, 'h2004f8, 'h100047, 'h1001e9, 'h1001ea, 'h1000ff, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1000fc, 'h1000fd, 'h1001f7, 'h10003c, 'h2004f8, 'h100047, 'h1000fe, 'h1001f8, 'h1000ff, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h1000fc, 'h10003c, 'h2004f8, 'h100047, 'h100207, 'h1000fd, 'h100208, 'h1000fe, 'h100209, 'h1000ff, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100213, 'h100214, 'h100215, 'h10003c, 'h2004f8, 'h100047, 'h100216, 'h1000fc, 'h100217, 'h1000fd, 'h100218, 'h1000fe, 'h100219, 'h1000ff, 'h10021a, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h10003c, 'h2004f8, 'h100047, 'h100227, 'h1000fc, 'h100228, 'h1000fd, 'h100229, 'h1000fe, 'h10022b, 'h1000ff, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h10003c, 'h2004f8, 'h100047, 'h100237, 'h1000fc, 'h100238, 'h1000fd, 'h100239, 'h1000fe, 'h10023a, 'h1000ff, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h10003c, 'h2004f8, 'h100047, 'h100245, 'h100246, 'h100247, 'h1000fc, 'h1000fd, 'h100248, 'h1000fe, 'h100249, 'h1000ff, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h10003c, 'h2004f8, 'h100047, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h1000fc, 'h1000fd, 'h100258, 'h1000fe, 'h100259, 'h1000ff, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h10003c, 'h2004f8, 'h100047, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h1000fc, 'h1000fd, 'h100268, 'h1000fe, 'h100269, 'h1000ff, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10003c, 'h2004f8, 'h100047, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h100103, 'h100100, 'h100101, 'h100172, 'h100102, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10003c, 'h2004f8, 'h100047, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100103, 'h100180, 'h100181, 'h100100, 'h100182, 'h100101, 'h100183, 'h100102, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h10003c, 'h2004f8, 'h100047, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h100103, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h100100, 'h100192, 'h100101, 'h100193, 'h100102, 'h100194, 'h100195, 'h100196, 'h10003c, 'h2004f8, 'h100047, 'h100197, 'h100198, 'h10019a, 'h10019b, 'h10019c, 'h100103, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h100100, 'h1001a3, 'h100101, 'h1001a4, 'h100102, 'h1001a6, 'h1001a7, 'h1001a8, 'h10003c, 'h2004f8, 'h100047, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h100103, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h100100, 'h100101, 'h1001b7, 'h100102, 'h1001b8, 'h10003c, 'h2004f8, 'h100047, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h100103, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h100100, 'h100101, 'h1001c7, 'h10003c, 'h2004f8, 'h100047, 'h100102, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h100103, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h100100, 'h10003c, 'h2004f8, 'h100047, 'h100101, 'h1001d7, 'h100102, 'h1001d8, 'h1001d9, 'h1001da, 'h100103, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h10003c, 'h2004f8, 'h100047, 'h1001e6, 'h100100, 'h100101, 'h1001e7, 'h100102, 'h1001e8, 'h100103, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h10003c, 'h2004f8, 'h100047, 'h1001f4, 'h1001f5, 'h1001f6, 'h100100, 'h100101, 'h1001f7, 'h100102, 'h1001f8, 'h100103, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h10003c, 'h2004f8, 'h100047, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100100, 'h100207, 'h100101, 'h100208, 'h100102, 'h100209, 'h100103, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h10003c, 'h2004f8, 'h100047, 'h100210, 'h100211, 'h100212, 'h100213, 'h100214, 'h100215, 'h100216, 'h100217, 'h100100, 'h100101, 'h100218, 'h100102, 'h100219, 'h100103, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h10003c, 'h2004f8, 'h100047, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h100100, 'h100101, 'h10022c, 'h100102, 'h10022d, 'h100103, 'h10022f, 'h100230, 'h100231, 'h10003c, 'h2004f8, 'h100047, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h100100, 'h100101, 'h10023c, 'h100102, 'h10023d, 'h100103, 'h10023e, 'h10023f, 'h10003c, 'h2004f8, 'h100047, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h100100, 'h100101, 'h10024c, 'h100102, 'h10024d, 'h100103, 'h10003c, 'h2004f8, 'h100047, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h100100, 'h100101, 'h10025c, 'h100102, 'h10003c, 'h2004f8, 'h100047, 'h10025d, 'h100103, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h100100, 'h100101, 'h10003c, 'h2004f8, 'h100047, 'h10026c, 'h100102, 'h10026d, 'h100103, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h100107, 'h100104, 'h100105, 'h100172, 'h100106, 'h100173, 'h100174, 'h100175, 'h10003c, 'h2004f8, 'h100047, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100107, 'h100180, 'h100181, 'h100104, 'h100105, 'h100182, 'h100106, 'h100183, 'h10003c, 'h2004f8, 'h100047, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h100107, 'h10018e, 'h10018f, 'h100190, 'h100191, 'h100192, 'h100104, 'h100105, 'h10003c, 'h2004f8, 'h100047, 'h100193, 'h100106, 'h100194, 'h100196, 'h100197, 'h100198, 'h10019a, 'h10019b, 'h10019c, 'h10019e, 'h100107, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h100104, 'h10003c, 'h2004f8, 'h100047, 'h100105, 'h1001a7, 'h100106, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h100107, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h100104, 'h10003c, 'h2004f8, 'h100047, 'h100105, 'h1001b7, 'h100106, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h100107, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h10003c, 'h2004f8, 'h100047, 'h1001c6, 'h100104, 'h100105, 'h1001c7, 'h100106, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h100107, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h10003c, 'h2004f8, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h100104, 'h100105, 'h1001d7, 'h100106, 'h1001d8, 'h1001d9, 'h1001da, 'h100107, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h10003c, 'h2004f8, 'h100047, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h100104, 'h100105, 'h1001e7, 'h100106, 'h1001e8, 'h100107, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h10003c, 'h2004f8, 'h100047, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h100104, 'h100105, 'h1001f7, 'h100106, 'h1001f8, 'h100107, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h10003c, 'h2004f8, 'h100047, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100104, 'h100207, 'h100105, 'h100208, 'h100106, 'h100209, 'h100107, 'h10020a, 'h10020b, 'h10003c, 'h2004f8, 'h100047, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100212, 'h100213, 'h100214, 'h100215, 'h100217, 'h100104, 'h100105, 'h100218, 'h100106, 'h100219, 'h100107, 'h10021b, 'h10003c, 'h2004f8, 'h100047, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h100104, 'h100105, 'h10022c, 'h100106, 'h10022d, 'h100107, 'h10003c, 'h2004f8, 'h100047, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h100104, 'h100105, 'h10023c, 'h100106, 'h10023d, 'h10003c, 'h2004f8, 'h100047, 'h100107, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h100104, 'h100105, 'h10024c, 'h10003c, 'h2004f8, 'h100047, 'h100106, 'h10024d, 'h100107, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h100104, 'h10003c, 'h2004f8, 'h100047, 'h100105, 'h10025c, 'h100106, 'h10025d, 'h100107, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10003c, 'h2004f8, 'h100047, 'h10026b, 'h100104, 'h100105, 'h10026c, 'h100106, 'h10026d, 'h100107, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h10010b, 'h100108, 'h100109, 'h100172, 'h10010a, 'h10003c, 'h2004f8, 'h100047, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h10010b, 'h100180, 'h100181, 'h100108, 'h100109, 'h10003c, 'h2004f8, 'h100047, 'h100182, 'h10010a, 'h100183, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018d, 'h10010b, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h10003c, 'h2004f8, 'h100047, 'h100108, 'h100109, 'h100193, 'h10010a, 'h100194, 'h100196, 'h100197, 'h100198, 'h10019a, 'h10019b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h10010b, 'h1001a2, 'h1001a3, 'h1001a4, 'h10003c, 'h2004f8, 'h100047, 'h1001a6, 'h100108, 'h100109, 'h1001a7, 'h10010a, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h10010b, 'h1001b3, 'h1001b4, 'h1001b5, 'h10003c, 'h2004f8, 'h100047, 'h1001b6, 'h100108, 'h100109, 'h1001b7, 'h10010a, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h10010b, 'h1001c1, 'h1001c2, 'h1001c3, 'h10003c, 'h2004f8, 'h100047, 'h1001c4, 'h1001c5, 'h1001c6, 'h100108, 'h100109, 'h1001c7, 'h10010a, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h10010b, 'h1001cf, 'h1001d0, 'h1001d1, 'h10003c, 'h2004f8, 'h100047, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h100108, 'h100109, 'h1001d7, 'h10010a, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h10010b, 'h1001dd, 'h1001de, 'h1001df, 'h10003c, 'h2004f8, 'h100047, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h100108, 'h100109, 'h1001e7, 'h10010a, 'h1001e8, 'h1001e9, 'h1001ea, 'h10010b, 'h1001eb, 'h1001ec, 'h1001ed, 'h10003c, 'h2004f8, 'h100047, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h100108, 'h100109, 'h1001f7, 'h10010a, 'h1001f8, 'h10010b, 'h1001f9, 'h1001fa, 'h1001fb, 'h10003c, 'h2004f8, 'h100047, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h100108, 'h100109, 'h100207, 'h10010a, 'h100208, 'h10010b, 'h100209, 'h10003c, 'h2004f8, 'h100047, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020e, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100108, 'h100109, 'h100218, 'h10010a, 'h100219, 'h10010b, 'h10003c, 'h2004f8, 'h100047, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h100108, 'h100109, 'h10022c, 'h10010a, 'h10022d, 'h10003c, 'h2004f8, 'h100047, 'h10010b, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h100108, 'h100109, 'h10023c, 'h10010a, 'h10003c, 'h2004f8, 'h100047, 'h10023d, 'h10010b, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h100108, 'h100109, 'h10003c, 'h2004f8, 'h100047, 'h10024c, 'h10010a, 'h10024d, 'h10010b, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10003c, 'h2004f8, 'h100047, 'h100108, 'h100109, 'h10025c, 'h10010a, 'h10025d, 'h10010b, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10003c, 'h2004f8, 'h100047, 'h10026a, 'h10026b, 'h100108, 'h100109, 'h10026c, 'h10010a, 'h10026d, 'h10010b, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h10010f, 'h10010d, 'h100172, 'h10010e, 'h10003c, 'h2004f8, 'h100047, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h10010f, 'h100181, 'h10010d, 'h100182, 'h10003c, 'h2004f8, 'h100047, 'h10010e, 'h100183, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h100189, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h10010f, 'h100192, 'h10010d, 'h100193, 'h10003c, 'h2004f8, 'h100047, 'h10010e, 'h100194, 'h100196, 'h100197, 'h100198, 'h10019a, 'h10019b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h10010f, 'h1001a6, 'h10010d, 'h1001a7, 'h10003c, 'h2004f8, 'h100047, 'h10010e, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h10010f, 'h1001b7, 'h10010d, 'h1001b8, 'h10003c, 'h2004f8, 'h100047, 'h10010e, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h10010f, 'h1001c6, 'h10010d, 'h1001c7, 'h10003c, 'h2004f8, 'h100047, 'h10010e, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h10010f, 'h1001d5, 'h1001d6, 'h10010d, 'h10003c, 'h2004f8, 'h100047, 'h1001d7, 'h10010e, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h10010f, 'h1001e5, 'h1001e6, 'h10003c, 'h2004f8, 'h100047, 'h10010d, 'h1001e7, 'h10010e, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h10010f, 'h1001f5, 'h10003c, 'h2004f8, 'h100047, 'h1001f6, 'h10010d, 'h1001f7, 'h10010e, 'h1001f8, 'h1001f9, 'h1001fa, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h10010f, 'h10003c, 'h2004f8, 'h100047, 'h100205, 'h100206, 'h10010d, 'h100207, 'h10010e, 'h100208, 'h100209, 'h10020a, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h10010f, 'h10003c, 'h2004f8, 'h100047, 'h100217, 'h100218, 'h10010d, 'h100219, 'h10010e, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10010f, 'h10003c, 'h2004f8, 'h100047, 'h10022b, 'h10022c, 'h10010d, 'h10022d, 'h10010e, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10010f, 'h10003c, 'h2004f8, 'h100047, 'h10023b, 'h10023c, 'h10010d, 'h10023d, 'h10010e, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10010f, 'h10003c, 'h2004f8, 'h100047, 'h10024a, 'h10024b, 'h10010d, 'h10024c, 'h10010e, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10003c, 'h2004f8, 'h100047, 'h10010f, 'h10025a, 'h10025b, 'h10010d, 'h10025c, 'h10010e, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h10003c, 'h2004f8, 'h100047, 'h100269, 'h10010f, 'h10026a, 'h10026b, 'h10010d, 'h10026c, 'h10010e, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100171, 'h100113, 'h100111, 'h100172, 'h100112, 'h10003c, 'h2004f8, 'h100047, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h100113, 'h100181, 'h100111, 'h100182, 'h10003c, 'h2004f8, 'h100047, 'h100112, 'h100183, 'h100184, 'h100185, 'h100186, 'h100187, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100113, 'h100193, 'h100194, 'h100196, 'h10003c, 'h2004f8, 'h100047, 'h100111, 'h100197, 'h100112, 'h100198, 'h10019a, 'h10019b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h100113, 'h1001a7, 'h1001a8, 'h1001aa, 'h10003c, 'h2004f8, 'h100047, 'h100111, 'h1001ab, 'h100112, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h100113, 'h1001b9, 'h1001ba, 'h10003c, 'h2004f8, 'h100047, 'h100111, 'h1001bb, 'h100112, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h100113, 'h1001c9, 'h10003c, 'h2004f8, 'h100047, 'h1001ca, 'h100111, 'h1001cb, 'h100112, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h100113, 'h10003c, 'h2004f8, 'h100047, 'h1001d9, 'h1001da, 'h100111, 'h1001db, 'h100112, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h10003c, 'h2004f8, 'h100047, 'h100113, 'h1001e9, 'h1001ea, 'h100111, 'h1001eb, 'h100112, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h10003c, 'h2004f8, 'h100047, 'h1001f8, 'h100113, 'h1001f9, 'h1001fa, 'h100111, 'h1001fb, 'h100112, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100206, 'h10003c, 'h2004f8, 'h100047, 'h100207, 'h100208, 'h100113, 'h100209, 'h10020b, 'h100111, 'h100112, 'h10020c, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10003c, 'h2004f8, 'h100047, 'h10021b, 'h10021c, 'h10021d, 'h100113, 'h10021f, 'h100111, 'h100220, 'h100112, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10003c, 'h2004f8, 'h100047, 'h10022f, 'h100230, 'h100231, 'h100113, 'h100232, 'h100233, 'h100111, 'h100234, 'h100112, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10003c, 'h2004f8, 'h100047, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100113, 'h100242, 'h100243, 'h100111, 'h100244, 'h100112, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10003c, 'h2004f8, 'h100047, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100113, 'h100252, 'h100253, 'h100111, 'h100254, 'h100112, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10003c, 'h2004f8, 'h100047, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100113, 'h100262, 'h100263, 'h100111, 'h100264, 'h100112, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10003c, 'h2004f8, 'h100047, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100113, 'h100272, 'h100171, 'h100117, 'h100115, 'h100172, 'h100116, 'h100173, 'h100174, 'h100175, 'h100176, 'h10003c, 'h2004f8, 'h100047, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h100117, 'h100181, 'h100182, 'h100115, 'h100116, 'h100183, 'h100184, 'h100186, 'h10003c, 'h2004f8, 'h100047, 'h100187, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100117, 'h100194, 'h100196, 'h100115, 'h100197, 'h100116, 'h100198, 'h10019a, 'h10003c, 'h2004f8, 'h100047, 'h10019b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h100117, 'h1001aa, 'h100115, 'h1001ab, 'h100116, 'h1001ac, 'h1001ae, 'h10003c, 'h2004f8, 'h100047, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h100117, 'h1001ba, 'h100115, 'h1001bb, 'h100116, 'h1001bc, 'h1001bd, 'h10003c, 'h2004f8, 'h100047, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h100117, 'h1001c9, 'h1001ca, 'h100115, 'h1001cb, 'h100116, 'h1001cc, 'h10003c, 'h2004f8, 'h100047, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h100117, 'h1001d9, 'h1001da, 'h100115, 'h1001db, 'h100116, 'h10003c, 'h2004f8, 'h100047, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h100117, 'h1001e9, 'h1001ea, 'h100115, 'h1001eb, 'h10003c, 'h2004f8, 'h100047, 'h100116, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h100117, 'h1001f9, 'h1001fa, 'h100115, 'h10003c, 'h2004f8, 'h100047, 'h1001fb, 'h100116, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h100201, 'h100202, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100117, 'h100209, 'h10020b, 'h100115, 'h10003c, 'h2004f8, 'h100047, 'h10020c, 'h100116, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h100117, 'h10021f, 'h100115, 'h10003c, 'h2004f8, 'h100047, 'h100220, 'h100116, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100117, 'h100232, 'h100233, 'h10003c, 'h2004f8, 'h100047, 'h100115, 'h100234, 'h100116, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100117, 'h100242, 'h10003c, 'h2004f8, 'h100047, 'h100243, 'h100115, 'h100244, 'h100116, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100117, 'h10003c, 'h2004f8, 'h100047, 'h100252, 'h100253, 'h100115, 'h100254, 'h100116, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h10003c, 'h2004f8, 'h100047, 'h100117, 'h100262, 'h100263, 'h100115, 'h100264, 'h100116, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h10003c, 'h2004f8, 'h100047, 'h100271, 'h100117, 'h100272, 'h100171, 'h10011b, 'h100119, 'h100172, 'h10011a, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10003c, 'h2004f8, 'h100047, 'h10017d, 'h10017e, 'h10017f, 'h100180, 'h10011b, 'h100182, 'h100119, 'h10011a, 'h100183, 'h100184, 'h100186, 'h100187, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h10003c, 'h2004f8, 'h100047, 'h100190, 'h100192, 'h100193, 'h100194, 'h10011b, 'h100196, 'h100119, 'h10011a, 'h100197, 'h100198, 'h10019a, 'h10019b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h10003c, 'h2004f8, 'h100047, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h10011b, 'h1001aa, 'h100119, 'h1001ab, 'h10011a, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h10003c, 'h2004f8, 'h100047, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h10011b, 'h1001ba, 'h100119, 'h1001bb, 'h10011a, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h10003c, 'h2004f8, 'h100047, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h10011b, 'h1001c9, 'h1001ca, 'h100119, 'h1001cb, 'h10011a, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h10003c, 'h2004f8, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h10011b, 'h1001d9, 'h1001da, 'h100119, 'h1001db, 'h10011a, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h10003c, 'h2004f8, 'h100047, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h10011b, 'h1001e9, 'h1001ea, 'h100119, 'h1001eb, 'h10011a, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h10003c, 'h2004f8, 'h100047, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h10011b, 'h1001f9, 'h1001fa, 'h100119, 'h1001fb, 'h10011a, 'h1001fc, 'h1001fd, 'h1001fe, 'h1001ff, 'h100200, 'h10003c, 'h2004f8, 'h100047, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h10011b, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h100119, 'h10011a, 'h100210, 'h100211, 'h100213, 'h100214, 'h10003c, 'h2004f8, 'h100047, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10011b, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100119, 'h100224, 'h10011a, 'h100225, 'h100227, 'h100228, 'h10003c, 'h2004f8, 'h100047, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h10011b, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100119, 'h100238, 'h10011a, 'h100239, 'h10003c, 'h2004f8, 'h100047, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h10011b, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100119, 'h100248, 'h10011a, 'h10003c, 'h2004f8, 'h100047, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h10011b, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100119, 'h100258, 'h10003c, 'h2004f8, 'h100047, 'h10011a, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h10011b, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100119, 'h10003c, 'h2004f8, 'h100047, 'h100268, 'h10011a, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h10011b, 'h100272, 'h100171, 'h10011f, 'h10011d, 'h100172, 'h10011e, 'h10003c, 'h2004f8, 'h100047, 'h100173, 'h100174, 'h100175, 'h100176, 'h100177, 'h100178, 'h100179, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h10011f, 'h10011d, 'h100183, 'h10011e, 'h10003c, 'h2004f8, 'h100047, 'h100184, 'h100186, 'h100187, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h10011f, 'h10011d, 'h100197, 'h10011e, 'h10003c, 'h2004f8, 'h100047, 'h100198, 'h10019a, 'h10019b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h10011f, 'h10011d, 'h1001ab, 'h10011e, 'h10003c, 'h2004f8, 'h100047, 'h1001ac, 'h1001ae, 'h1001af, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h10011f, 'h10011d, 'h1001bb, 'h10011e, 'h10003c, 'h2004f8, 'h100047, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h10011f, 'h1001ca, 'h10011d, 'h1001cb, 'h10003c, 'h2004f8, 'h100047, 'h10011e, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h10011f, 'h1001d9, 'h1001da, 'h10011d, 'h10003c, 'h2004f8, 'h100047, 'h1001db, 'h10011e, 'h1001dc, 'h1001dd, 'h1001de, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h10011f, 'h1001e9, 'h1001ea, 'h10003c, 'h2004f8, 'h100047, 'h10011d, 'h1001eb, 'h10011e, 'h1001ec, 'h1001ed, 'h1001ee, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f6, 'h1001f7, 'h1001f8, 'h10011f, 'h1001f9, 'h10003c, 'h2004f8, 'h100047, 'h1001fa, 'h1001fb, 'h10011d, 'h10011e, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10011f, 'h10020c, 'h10003c, 'h2004f8, 'h100047, 'h10020d, 'h10020f, 'h10011d, 'h10011e, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h10011f, 'h100220, 'h10003c, 'h2004f8, 'h100047, 'h100221, 'h100223, 'h10011d, 'h100224, 'h10011e, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h10011f, 'h100233, 'h10003c, 'h2004f8, 'h100047, 'h100234, 'h100235, 'h100236, 'h100237, 'h10011d, 'h100238, 'h10011e, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h10011f, 'h100242, 'h10003c, 'h2004f8, 'h100047, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h10011d, 'h100248, 'h10011e, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h10011f, 'h10003c, 'h2004f8, 'h100047, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h10011d, 'h100258, 'h10011e, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h10003c, 'h2004f8, 'h100047, 'h10011f, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h10011d, 'h100268, 'h10011e, 'h100269, 'h10026a, 'h10026b, 'h10026c, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h10003c, 'h2004f8, 'h100047, 'h100271, 'h10011f, 'h100272, 'h100171, 'h100123, 'h100173, 'h100121, 'h100172, 'h100122, 'h100174, 'h100175, 'h100177, 'h100176, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h10003c, 'h2004f8, 'h100047, 'h100180, 'h100182, 'h100183, 'h100123, 'h100184, 'h100186, 'h100187, 'h100121, 'h100122, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100194, 'h10003c, 'h2004f8, 'h100047, 'h100193, 'h100196, 'h100198, 'h100123, 'h100197, 'h10019a, 'h10019c, 'h100121, 'h100122, 'h10019b, 'h10019e, 'h1001a0, 'h10019f, 'h1001a2, 'h1001a4, 'h1001a3, 'h1001a6, 'h1001a8, 'h10003c, 'h2004f8, 'h100047, 'h1001a7, 'h1001aa, 'h1001ac, 'h100123, 'h1001ab, 'h1001ae, 'h1001b0, 'h100121, 'h1001af, 'h100122, 'h1001b1, 'h1001b2, 'h1001b4, 'h1001b3, 'h1001b5, 'h1001b6, 'h1001b8, 'h1001b7, 'h10003c, 'h2004f8, 'h100047, 'h1001b9, 'h1001ba, 'h1001bc, 'h100123, 'h1001bb, 'h1001bd, 'h1001be, 'h1001c0, 'h100121, 'h1001bf, 'h100122, 'h1001c1, 'h1001c2, 'h1001c4, 'h1001c3, 'h1001c5, 'h1001c6, 'h1001c8, 'h10003c, 'h2004f8, 'h100047, 'h1001c7, 'h1001c9, 'h1001ca, 'h100123, 'h1001cc, 'h1001cb, 'h1001cd, 'h1001ce, 'h1001d0, 'h100121, 'h1001cf, 'h100122, 'h1001d1, 'h1001d2, 'h1001d4, 'h1001d3, 'h1001d5, 'h1001d6, 'h1001d8, 'h10003c, 'h2004f8, 'h100047, 'h1001d7, 'h1001d9, 'h100123, 'h1001da, 'h1001dc, 'h1001db, 'h1001dd, 'h1001de, 'h1001e0, 'h100121, 'h1001df, 'h100122, 'h1001e1, 'h1001e2, 'h1001e4, 'h1001e3, 'h1001e5, 'h1001e6, 'h1001e8, 'h10003c, 'h2004f8, 'h100047, 'h1001e7, 'h100123, 'h1001e9, 'h1001ea, 'h1001ec, 'h1001eb, 'h1001ed, 'h1001ee, 'h1001f0, 'h100121, 'h1001ef, 'h100122, 'h1001f1, 'h1001f2, 'h1001f4, 'h1001f3, 'h1001f5, 'h1001f6, 'h1001f8, 'h10003c, 'h2004f8, 'h100047, 'h100123, 'h1001f7, 'h1001f9, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h100121, 'h100201, 'h100203, 'h100204, 'h100122, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h10003c, 'h2004f8, 'h100047, 'h100123, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100215, 'h100121, 'h100214, 'h100217, 'h100219, 'h100122, 'h100218, 'h10021b, 'h10021d, 'h10021c, 'h10021f, 'h100221, 'h10003c, 'h2004f8, 'h100047, 'h100123, 'h100220, 'h100223, 'h100225, 'h100224, 'h100227, 'h100229, 'h100121, 'h100228, 'h10022b, 'h10022d, 'h10022c, 'h100122, 'h10022f, 'h100231, 'h100230, 'h100232, 'h100233, 'h100235, 'h10003c, 'h2004f8, 'h100047, 'h100123, 'h100234, 'h100236, 'h100237, 'h100239, 'h100238, 'h100121, 'h10023a, 'h10023b, 'h10023d, 'h10023c, 'h100122, 'h10023e, 'h10023f, 'h100241, 'h100240, 'h100242, 'h100243, 'h100245, 'h10003c, 'h2004f8, 'h100047, 'h100123, 'h100244, 'h100246, 'h100247, 'h100249, 'h100121, 'h100248, 'h10024a, 'h10024b, 'h10024d, 'h10024c, 'h100122, 'h10024e, 'h10024f, 'h100251, 'h100250, 'h100252, 'h100253, 'h100255, 'h10003c, 'h2004f8, 'h100047, 'h100123, 'h100254, 'h100256, 'h100257, 'h100259, 'h100121, 'h100258, 'h10025a, 'h10025b, 'h10025d, 'h10025c, 'h100122, 'h10025e, 'h10025f, 'h100261, 'h100260, 'h100262, 'h100263, 'h100265, 'h10003c, 'h2004f8, 'h100047, 'h100123, 'h100264, 'h100266, 'h100267, 'h100269, 'h100121, 'h100268, 'h10026a, 'h10026b, 'h10026d, 'h10026c, 'h100122, 'h10026e, 'h10026f, 'h100271, 'h100270, 'h100272, 'h100171, 'h100127, 'h10003c, 'h2004f8, 'h100047, 'h100172, 'h100125, 'h100126, 'h100173, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100127, 'h10003c, 'h2004f8, 'h100047, 'h100186, 'h100125, 'h100126, 'h100187, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h100127, 'h10003c, 'h2004f8, 'h100047, 'h10019a, 'h100125, 'h100126, 'h10019b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h100127, 'h10003c, 'h2004f8, 'h100047, 'h1001ae, 'h100125, 'h1001af, 'h100126, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h100127, 'h10003c, 'h2004f8, 'h100047, 'h1001bd, 'h1001be, 'h100125, 'h1001bf, 'h100126, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h10003c, 'h2004f8, 'h100047, 'h100127, 'h1001cd, 'h1001ce, 'h100125, 'h1001cf, 'h100126, 'h1001d0, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h10003c, 'h2004f8, 'h100047, 'h1001dc, 'h100127, 'h1001dd, 'h1001de, 'h100125, 'h1001df, 'h100126, 'h1001e0, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h10003c, 'h2004f8, 'h100047, 'h1001eb, 'h1001ec, 'h100127, 'h1001ed, 'h1001ee, 'h100125, 'h1001ef, 'h100126, 'h1001f0, 'h1001f1, 'h1001f2, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fb, 'h10003c, 'h2004f8, 'h100047, 'h1001fc, 'h1001fd, 'h100127, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100125, 'h100126, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h10003c, 'h2004f8, 'h100047, 'h100210, 'h100211, 'h100127, 'h100213, 'h100214, 'h100215, 'h100217, 'h100125, 'h100126, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h10003c, 'h2004f8, 'h100047, 'h100224, 'h100225, 'h100127, 'h100227, 'h100228, 'h100229, 'h10022b, 'h100125, 'h10022c, 'h100126, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h10003c, 'h2004f8, 'h100047, 'h100236, 'h100237, 'h100127, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h100125, 'h10023c, 'h100126, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h10003c, 'h2004f8, 'h100047, 'h100245, 'h100246, 'h100127, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h100125, 'h10024c, 'h100126, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h10003c, 'h2004f8, 'h100047, 'h100254, 'h100255, 'h100127, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h100125, 'h10025c, 'h100126, 'h10025d, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h10003c, 'h2004f8, 'h100047, 'h100263, 'h100264, 'h100265, 'h100127, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h100125, 'h10026c, 'h100126, 'h10026d, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h10003c, 'h2004f8, 'h100047, 'h100272, 'h100172, 'h10012c, 'h100129, 'h10012a, 'h100173, 'h10012b, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h10003c, 'h2004f8, 'h100047, 'h100183, 'h100184, 'h100186, 'h10012c, 'h100129, 'h10012a, 'h100187, 'h10012b, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h10003c, 'h2004f8, 'h100047, 'h100196, 'h100197, 'h100198, 'h10019a, 'h10012c, 'h100129, 'h10012a, 'h10019b, 'h10012b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h10003c, 'h2004f8, 'h100047, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h10012c, 'h100129, 'h1001af, 'h10012a, 'h1001b0, 'h10012b, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h2004f8, 'h100047, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h10012c, 'h100129, 'h1001bf, 'h10012a, 'h1001c0, 'h10012b, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h10003c, 'h2004f8, 'h100047, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h10012c, 'h100129, 'h1001cf, 'h10012a, 'h1001d0, 'h10012b, 'h1001d1, 'h1001d2, 'h1001d3, 'h10003c, 'h2004f8, 'h100047, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001de, 'h10012c, 'h100129, 'h1001df, 'h10012a, 'h1001e0, 'h10012b, 'h1001e1, 'h10003c, 'h2004f8, 'h100047, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ee, 'h10012c, 'h1001ef, 'h100129, 'h10012a, 'h1001f0, 'h10003c, 'h2004f8, 'h100047, 'h10012b, 'h1001f1, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h10012c, 'h100129, 'h10012a, 'h10003c, 'h2004f8, 'h100047, 'h100204, 'h10012b, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h10012c, 'h100129, 'h10003c, 'h2004f8, 'h100047, 'h10012a, 'h100218, 'h10012b, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10012c, 'h10003c, 'h2004f8, 'h100047, 'h100129, 'h10022c, 'h10012a, 'h10022d, 'h10012b, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10012c, 'h10003c, 'h2004f8, 'h100047, 'h100129, 'h10023c, 'h10012a, 'h10023d, 'h10012b, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10003c, 'h2004f8, 'h100047, 'h10024b, 'h10012c, 'h100129, 'h10024c, 'h10012a, 'h10024d, 'h10012b, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h10003c, 'h2004f8, 'h100047, 'h100259, 'h10025a, 'h10025b, 'h10012c, 'h100129, 'h10025c, 'h10012a, 'h10025d, 'h10012b, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h10003c, 'h2004f8, 'h100047, 'h100267, 'h100268, 'h100269, 'h10026a, 'h10026b, 'h10012c, 'h100129, 'h10026c, 'h10012a, 'h10026d, 'h10012b, 'h10026e, 'h10026f, 'h100270, 'h100271, 'h100272, 'h100172, 'h100130, 'h10003c, 'h2004f8, 'h100047, 'h10012d, 'h10012e, 'h100173, 'h10012f, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100130, 'h10003c, 'h2004f8, 'h100047, 'h100186, 'h10012d, 'h10012e, 'h100187, 'h10012f, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h10003c, 'h2004f8, 'h100047, 'h100130, 'h10019a, 'h10012d, 'h10012e, 'h10019b, 'h10012f, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h10003c, 'h2004f8, 'h100047, 'h1001ac, 'h100130, 'h1001ae, 'h10012d, 'h1001af, 'h10012e, 'h1001b0, 'h10012f, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h10003c, 'h2004f8, 'h100047, 'h1001bb, 'h1001bc, 'h1001bd, 'h100130, 'h1001be, 'h10012d, 'h1001bf, 'h10012e, 'h1001c0, 'h10012f, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h10003c, 'h2004f8, 'h100047, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h100130, 'h1001ce, 'h10012d, 'h1001cf, 'h10012e, 'h1001d0, 'h10012f, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h10003c, 'h2004f8, 'h100047, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h100130, 'h1001de, 'h10012d, 'h1001df, 'h10012e, 'h1001e0, 'h10012f, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h10003c, 'h2004f8, 'h100047, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001ea, 'h1001eb, 'h1001ec, 'h1001ed, 'h100130, 'h1001ef, 'h10012d, 'h10012e, 'h1001f0, 'h10012f, 'h1001f1, 'h1001f3, 'h1001f4, 'h10003c, 'h2004f8, 'h100047, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100130, 'h100203, 'h10012d, 'h10012e, 'h100204, 'h10012f, 'h100205, 'h100207, 'h10003c, 'h2004f8, 'h100047, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100130, 'h100217, 'h10012d, 'h10012e, 'h100218, 'h10012f, 'h100219, 'h10003c, 'h2004f8, 'h100047, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h100130, 'h10022b, 'h10012d, 'h10012e, 'h10022c, 'h10012f, 'h10003c, 'h2004f8, 'h100047, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h100130, 'h10023b, 'h10012d, 'h10023c, 'h10012e, 'h10003c, 'h2004f8, 'h100047, 'h10023d, 'h10012f, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h100130, 'h10024b, 'h10012d, 'h10003c, 'h2004f8, 'h100047, 'h10024c, 'h10012e, 'h10024d, 'h10012f, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h100130, 'h10003c, 'h2004f8, 'h100047, 'h10025b, 'h10012d, 'h10025c, 'h10012e, 'h10025d, 'h10012f, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10003c, 'h2004f8, 'h100047, 'h10026a, 'h100130, 'h10026b, 'h10026c, 'h10012d, 'h10012e, 'h10026d, 'h10012f, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100134, 'h100131, 'h100132, 'h100173, 'h100133, 'h10003c, 'h2004f8, 'h100047, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100134, 'h100186, 'h100131, 'h100132, 'h100187, 'h10003c, 'h2004f8, 'h100047, 'h100133, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h100134, 'h10019a, 'h100131, 'h100132, 'h10003c, 'h2004f8, 'h100047, 'h10019b, 'h100133, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h100134, 'h1001ae, 'h100131, 'h10003c, 'h2004f8, 'h100047, 'h100132, 'h1001af, 'h100133, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h100134, 'h10003c, 'h2004f8, 'h100047, 'h1001be, 'h100131, 'h1001bf, 'h100132, 'h1001c0, 'h100133, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h10003c, 'h2004f8, 'h100047, 'h1001cd, 'h100134, 'h1001ce, 'h100131, 'h1001cf, 'h100132, 'h1001d0, 'h100133, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h10003c, 'h2004f8, 'h100047, 'h1001db, 'h1001dc, 'h1001dd, 'h100134, 'h1001de, 'h100131, 'h1001df, 'h100132, 'h1001e0, 'h100133, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e6, 'h1001e7, 'h1001e8, 'h10003c, 'h2004f8, 'h100047, 'h1001e9, 'h1001eb, 'h1001ec, 'h1001ed, 'h100134, 'h1001ef, 'h100131, 'h100132, 'h1001f0, 'h100133, 'h1001f1, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fb, 'h10003c, 'h2004f8, 'h100047, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100134, 'h100203, 'h100131, 'h100132, 'h100204, 'h100133, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h10020d, 'h10003c, 'h2004f8, 'h100047, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100134, 'h100217, 'h100131, 'h100132, 'h100218, 'h100133, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h10003c, 'h2004f8, 'h100047, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h100134, 'h10022b, 'h100131, 'h100132, 'h10022c, 'h100133, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h10003c, 'h2004f8, 'h100047, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h100134, 'h10023b, 'h100131, 'h10023c, 'h100132, 'h10023d, 'h100133, 'h10023e, 'h10023f, 'h100240, 'h10003c, 'h2004f8, 'h100047, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h100134, 'h10024b, 'h100131, 'h10024c, 'h100132, 'h10024d, 'h100133, 'h10024e, 'h10003c, 'h2004f8, 'h100047, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h100134, 'h10025b, 'h100131, 'h10025c, 'h100132, 'h10025d, 'h10003c, 'h2004f8, 'h100047, 'h100133, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h100264, 'h100265, 'h100266, 'h100267, 'h100268, 'h100269, 'h10026a, 'h100134, 'h10026c, 'h100131, 'h100132, 'h10003c, 'h2004f8, 'h100047, 'h10026d, 'h100133, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100138, 'h100135, 'h100136, 'h100173, 'h100137, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10003c, 'h2004f8, 'h100047, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100138, 'h100186, 'h100135, 'h100136, 'h100187, 'h100137, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10003c, 'h2004f8, 'h100047, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h100138, 'h10019a, 'h100135, 'h100136, 'h10019b, 'h100137, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h10003c, 'h2004f8, 'h100047, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h100138, 'h1001ae, 'h100135, 'h100136, 'h1001af, 'h100137, 'h1001b0, 'h1001b1, 'h1001b2, 'h10003c, 'h2004f8, 'h100047, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h100138, 'h1001be, 'h100135, 'h1001bf, 'h100136, 'h1001c0, 'h100137, 'h10003c, 'h2004f8, 'h100047, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h100138, 'h1001ce, 'h100135, 'h1001cf, 'h100136, 'h10003c, 'h2004f8, 'h100047, 'h1001d0, 'h100137, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h100138, 'h1001de, 'h100135, 'h10003c, 'h2004f8, 'h100047, 'h1001df, 'h100136, 'h1001e0, 'h100137, 'h1001e1, 'h1001e2, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001eb, 'h1001ec, 'h1001ed, 'h100138, 'h1001ef, 'h100135, 'h10003c, 'h2004f8, 'h100047, 'h1001f0, 'h100136, 'h1001f1, 'h100137, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100138, 'h100203, 'h10003c, 'h2004f8, 'h100047, 'h100135, 'h100136, 'h100204, 'h100137, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100138, 'h10003c, 'h2004f8, 'h100047, 'h100217, 'h100135, 'h100136, 'h100218, 'h100137, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10003c, 'h2004f8, 'h100047, 'h100138, 'h10022b, 'h100135, 'h100136, 'h10022c, 'h100137, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10003c, 'h2004f8, 'h100047, 'h10023a, 'h100138, 'h10023b, 'h100135, 'h10023c, 'h100136, 'h10023d, 'h100137, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100247, 'h10003c, 'h2004f8, 'h100047, 'h100248, 'h100249, 'h10024a, 'h100138, 'h10024b, 'h100135, 'h10024c, 'h100136, 'h10024d, 'h100137, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100255, 'h10003c, 'h2004f8, 'h100047, 'h100256, 'h100257, 'h100258, 'h100259, 'h10025a, 'h100138, 'h10025b, 'h100135, 'h10025c, 'h100136, 'h10025d, 'h100137, 'h10025e, 'h10025f, 'h100260, 'h100261, 'h100262, 'h100263, 'h10003c, 'h2004f8, 'h100047, 'h100264, 'h100265, 'h100266, 'h100268, 'h100269, 'h10026a, 'h100138, 'h10026c, 'h100135, 'h100136, 'h10026d, 'h100137, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h10013c, 'h100173, 'h10003c, 'h2004f8, 'h100047, 'h100139, 'h10013a, 'h10013b, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h10013c, 'h100186, 'h100187, 'h10003c, 'h2004f8, 'h100047, 'h100139, 'h10013a, 'h10013b, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h10013c, 'h100198, 'h10019a, 'h10019b, 'h10003c, 'h2004f8, 'h100047, 'h100139, 'h10013a, 'h10013b, 'h10019c, 'h10019e, 'h1001a0, 'h10019f, 'h1001a2, 'h1001a4, 'h1001a3, 'h1001a6, 'h1001a8, 'h1001a7, 'h1001aa, 'h10013c, 'h1001ac, 'h1001ab, 'h1001ae, 'h1001b0, 'h10003c, 'h2004f8, 'h100047, 'h100139, 'h10013a, 'h1001af, 'h10013b, 'h1001b1, 'h1001b2, 'h1001b4, 'h1001b3, 'h1001b5, 'h1001b6, 'h1001b8, 'h1001b7, 'h1001b9, 'h10013c, 'h1001ba, 'h1001bc, 'h1001bb, 'h1001bd, 'h10003c, 'h2004f8, 'h100047, 'h1001be, 'h1001c0, 'h100139, 'h1001bf, 'h10013a, 'h10013b, 'h1001c1, 'h1001c2, 'h1001c4, 'h1001c3, 'h1001c5, 'h1001c6, 'h1001c8, 'h10013c, 'h1001c7, 'h1001c9, 'h1001ca, 'h1001cc, 'h10003c, 'h2004f8, 'h100047, 'h1001cb, 'h1001cd, 'h1001ce, 'h1001d0, 'h100139, 'h1001cf, 'h10013a, 'h10013b, 'h1001d1, 'h1001d2, 'h1001d4, 'h1001d3, 'h1001d5, 'h10013c, 'h1001d6, 'h1001d8, 'h1001d7, 'h1001d9, 'h10003c, 'h2004f8, 'h100047, 'h1001da, 'h1001dc, 'h1001db, 'h1001dd, 'h1001de, 'h1001e0, 'h1001df, 'h100139, 'h10013a, 'h10013b, 'h1001e1, 'h1001e3, 'h1001e4, 'h10013c, 'h1001e5, 'h1001e7, 'h1001e8, 'h1001e9, 'h10003c, 'h2004f8, 'h100047, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h100139, 'h10013a, 'h10013b, 'h1001f5, 'h1001f7, 'h10013c, 'h1001f8, 'h1001f9, 'h1001fb, 'h1001fc, 'h10003c, 'h2004f8, 'h100047, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100139, 'h10013a, 'h10013b, 'h100209, 'h10013c, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h100210, 'h10003c, 'h2004f8, 'h100047, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h100139, 'h10013a, 'h10013b, 'h10021d, 'h10013c, 'h10021f, 'h100221, 'h100220, 'h100223, 'h100225, 'h10003c, 'h2004f8, 'h100047, 'h100224, 'h100227, 'h100229, 'h100228, 'h10022b, 'h10022d, 'h10022c, 'h10022f, 'h100231, 'h100139, 'h10013a, 'h100230, 'h10013b, 'h10013c, 'h100232, 'h100233, 'h100235, 'h100234, 'h10003c, 'h2004f8, 'h100047, 'h100236, 'h100237, 'h100239, 'h100238, 'h10023a, 'h10023b, 'h10023d, 'h10023c, 'h10023e, 'h10023f, 'h100241, 'h100139, 'h100240, 'h10013a, 'h10013b, 'h100242, 'h10013c, 'h100243, 'h100245, 'h10003c, 'h2004f8, 'h100047, 'h100244, 'h100246, 'h100247, 'h100249, 'h100248, 'h10024a, 'h10024b, 'h10024d, 'h10024c, 'h10024e, 'h10024f, 'h100251, 'h100139, 'h100250, 'h10013a, 'h10013b, 'h100252, 'h10013c, 'h10003c, 'h2004f8, 'h100047, 'h100253, 'h100255, 'h100254, 'h100256, 'h100257, 'h100259, 'h100258, 'h10025a, 'h10025b, 'h10025d, 'h10025c, 'h10025e, 'h10025f, 'h100261, 'h100260, 'h100139, 'h10013a, 'h10013b, 'h10003c, 'h2004f8, 'h100047, 'h100262, 'h10013c, 'h100264, 'h100265, 'h100266, 'h100268, 'h100269, 'h10026a, 'h10026c, 'h10026d, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100140, 'h10013d, 'h10013e, 'h10003c, 'h2004f8, 'h100047, 'h100173, 'h10013f, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100140, 'h100186, 'h10013d, 'h10003c, 'h2004f8, 'h100047, 'h10013e, 'h100187, 'h10013f, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h100140, 'h10019a, 'h10003c, 'h2004f8, 'h100047, 'h10013d, 'h10013e, 'h10019b, 'h10013f, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h100140, 'h10003c, 'h2004f8, 'h100047, 'h1001ae, 'h10013d, 'h10013e, 'h1001af, 'h10013f, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h10003c, 'h2004f8, 'h100047, 'h100140, 'h1001bd, 'h1001be, 'h10013d, 'h1001bf, 'h10013e, 'h1001c0, 'h10013f, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h10003c, 'h2004f8, 'h100047, 'h100140, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h10013d, 'h1001cf, 'h10013e, 'h1001d0, 'h10013f, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d6, 'h1001d7, 'h1001d8, 'h10003c, 'h2004f8, 'h100047, 'h1001d9, 'h100140, 'h1001da, 'h1001db, 'h1001dc, 'h1001dd, 'h1001df, 'h10013d, 'h10013e, 'h1001e0, 'h10013f, 'h1001e1, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e7, 'h1001e8, 'h1001e9, 'h10003c, 'h2004f8, 'h100047, 'h1001eb, 'h100140, 'h1001ec, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h10013d, 'h10013e, 'h1001f4, 'h10013f, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h1001fb, 'h1001fc, 'h10003c, 'h2004f8, 'h100047, 'h1001fd, 'h100140, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h10013d, 'h10013e, 'h100208, 'h10013f, 'h100209, 'h10020b, 'h10020c, 'h10020d, 'h10020f, 'h10003c, 'h2004f8, 'h100047, 'h100210, 'h100211, 'h100140, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10013d, 'h10013e, 'h10021c, 'h10013f, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h10003c, 'h2004f8, 'h100047, 'h100223, 'h100224, 'h100225, 'h100140, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h10013d, 'h10013e, 'h100230, 'h10013f, 'h100231, 'h100232, 'h100233, 'h10003c, 'h2004f8, 'h100047, 'h100234, 'h100235, 'h100236, 'h100140, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h10013d, 'h100240, 'h10013e, 'h100241, 'h10013f, 'h10003c, 'h2004f8, 'h100047, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100140, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h10024f, 'h10013d, 'h100250, 'h10013e, 'h10003c, 'h2004f8, 'h100047, 'h100251, 'h10013f, 'h100252, 'h100253, 'h100254, 'h100255, 'h100256, 'h100140, 'h100257, 'h100258, 'h100259, 'h10025a, 'h10025b, 'h10025c, 'h10025d, 'h10025e, 'h100260, 'h10013d, 'h10003c, 'h2004f8, 'h100047, 'h10013e, 'h100261, 'h10013f, 'h100262, 'h100264, 'h100265, 'h100266, 'h100140, 'h100268, 'h100269, 'h10026a, 'h10026c, 'h10026d, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100144, 'h100173, 'h10003c, 'h2004f8, 'h100047, 'h100141, 'h100142, 'h100143, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100144, 'h100186, 'h100187, 'h10003c, 'h2004f8, 'h100047, 'h100141, 'h100142, 'h100143, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100144, 'h100198, 'h10019a, 'h10019b, 'h10003c, 'h2004f8, 'h100047, 'h100141, 'h100142, 'h100143, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a8, 'h1001a7, 'h1001aa, 'h100144, 'h1001ac, 'h1001ab, 'h1001ae, 'h1001b0, 'h10003c, 'h2004f8, 'h100047, 'h100141, 'h100142, 'h1001af, 'h100143, 'h1001b1, 'h1001b2, 'h1001b4, 'h1001b3, 'h1001b5, 'h1001b6, 'h1001b8, 'h1001b7, 'h1001b9, 'h100144, 'h1001ba, 'h1001bc, 'h1001bb, 'h1001bd, 'h10003c, 'h2004f8, 'h100047, 'h1001be, 'h1001c0, 'h100141, 'h100142, 'h1001bf, 'h100143, 'h1001c1, 'h1001c2, 'h1001c4, 'h1001c3, 'h1001c5, 'h1001c6, 'h1001c8, 'h100144, 'h1001c7, 'h1001c9, 'h1001ca, 'h1001cc, 'h10003c, 'h2004f8, 'h100047, 'h1001cb, 'h1001cd, 'h1001ce, 'h1001d0, 'h100141, 'h1001cf, 'h100142, 'h100143, 'h1001d1, 'h1001d2, 'h1001d4, 'h1001d3, 'h1001d5, 'h100144, 'h1001d6, 'h1001d8, 'h1001d7, 'h1001d9, 'h10003c, 'h2004f8, 'h100047, 'h1001db, 'h1001dc, 'h1001dd, 'h1001df, 'h1001e0, 'h100141, 'h100142, 'h100143, 'h1001e1, 'h1001e3, 'h1001e4, 'h1001e5, 'h1001e7, 'h100144, 'h1001e8, 'h1001e9, 'h1001eb, 'h1001ec, 'h10003c, 'h2004f8, 'h100047, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h100141, 'h100142, 'h100143, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h100144, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h10003c, 'h2004f8, 'h100047, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100141, 'h100142, 'h100143, 'h100209, 'h10020b, 'h10020c, 'h100144, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h10003c, 'h2004f8, 'h100047, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h100141, 'h100142, 'h100143, 'h10021d, 'h10021f, 'h100144, 'h100220, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100229, 'h10003c, 'h2004f8, 'h100047, 'h100228, 'h10022b, 'h10022d, 'h10022c, 'h10022f, 'h100231, 'h100141, 'h100142, 'h100230, 'h100143, 'h100144, 'h100232, 'h100233, 'h100235, 'h100234, 'h100236, 'h100237, 'h100239, 'h10003c, 'h2004f8, 'h100047, 'h100238, 'h10023a, 'h10023b, 'h10023d, 'h10023c, 'h10023e, 'h10023f, 'h100241, 'h100141, 'h100142, 'h100240, 'h100143, 'h100144, 'h100242, 'h100243, 'h100245, 'h100244, 'h100246, 'h10003c, 'h2004f8, 'h100047, 'h100247, 'h100249, 'h100248, 'h10024a, 'h10024b, 'h10024d, 'h10024c, 'h10024e, 'h10024f, 'h100251, 'h100141, 'h100250, 'h100142, 'h100143, 'h100252, 'h100144, 'h100253, 'h100255, 'h10003c, 'h2004f8, 'h100047, 'h100254, 'h100256, 'h100257, 'h100259, 'h100258, 'h10025a, 'h10025c, 'h10025d, 'h10025e, 'h100260, 'h100261, 'h100141, 'h100142, 'h100143, 'h100262, 'h100144, 'h100264, 'h100265, 'h10003c, 'h2004f8, 'h100047, 'h100266, 'h100268, 'h100269, 'h10026a, 'h10026c, 'h10026d, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100148, 'h100173, 'h100145, 'h100146, 'h100147, 'h100174, 'h100176, 'h100177, 'h10003c, 'h2004f8, 'h100047, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100148, 'h100186, 'h100187, 'h100145, 'h100146, 'h100147, 'h100188, 'h10018a, 'h10018b, 'h10003c, 'h2004f8, 'h100047, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100148, 'h100198, 'h10019a, 'h10019b, 'h100145, 'h100146, 'h100147, 'h10019c, 'h10019e, 'h10019f, 'h10003c, 'h2004f8, 'h100047, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h100148, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h100145, 'h100146, 'h100147, 'h1001b0, 'h1001b1, 'h10003c, 'h2004f8, 'h100047, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h100148, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h1001be, 'h1001bf, 'h100145, 'h100146, 'h100147, 'h10003c, 'h2004f8, 'h100047, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h100148, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001ce, 'h1001cf, 'h100145, 'h10003c, 'h2004f8, 'h100047, 'h100146, 'h1001d0, 'h100147, 'h1001d1, 'h1001d2, 'h1001d3, 'h1001d4, 'h1001d5, 'h100148, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001db, 'h1001dc, 'h1001dd, 'h1001df, 'h1001e0, 'h1001e1, 'h10003c, 'h2004f8, 'h100047, 'h1001e3, 'h100145, 'h100146, 'h1001e4, 'h100147, 'h1001e5, 'h1001e7, 'h1001e8, 'h1001e9, 'h100148, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h10003c, 'h2004f8, 'h100047, 'h1001f5, 'h1001f7, 'h1001f8, 'h100145, 'h100146, 'h100147, 'h1001f9, 'h1001fb, 'h1001fc, 'h100148, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h10003c, 'h2004f8, 'h100047, 'h100209, 'h10020b, 'h10020c, 'h100145, 'h100146, 'h100147, 'h10020d, 'h10020f, 'h100148, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10003c, 'h2004f8, 'h100047, 'h10021d, 'h10021f, 'h100220, 'h100145, 'h100146, 'h100147, 'h100221, 'h100148, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h10003c, 'h2004f8, 'h100047, 'h100231, 'h100232, 'h100233, 'h100234, 'h100145, 'h100146, 'h100147, 'h100235, 'h100148, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10003c, 'h2004f8, 'h100047, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100243, 'h100244, 'h100145, 'h100146, 'h100147, 'h100245, 'h100148, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10003c, 'h2004f8, 'h100047, 'h10024d, 'h10024e, 'h10024f, 'h100250, 'h100251, 'h100252, 'h100253, 'h100254, 'h100145, 'h100146, 'h100255, 'h100147, 'h100256, 'h100148, 'h100258, 'h100259, 'h10025a, 'h10025c, 'h10003c, 'h2004f8, 'h100047, 'h10025d, 'h10025e, 'h100260, 'h100261, 'h100262, 'h100264, 'h100265, 'h100266, 'h100268, 'h100145, 'h100146, 'h100269, 'h100147, 'h10026a, 'h100148, 'h10026c, 'h10026d, 'h10026e, 'h10003c, 'h2004f8, 'h100047, 'h100270, 'h100271, 'h100272, 'h100172, 'h10014c, 'h100173, 'h100149, 'h10014a, 'h10014b, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h10003c, 'h2004f8, 'h100047, 'h100180, 'h100182, 'h100183, 'h100184, 'h10014c, 'h100186, 'h100187, 'h100149, 'h10014a, 'h10014b, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h10003c, 'h2004f8, 'h100047, 'h100194, 'h100196, 'h100197, 'h10014c, 'h100198, 'h10019a, 'h10019b, 'h100149, 'h10014a, 'h10014b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h10003c, 'h2004f8, 'h100047, 'h1001a8, 'h1001aa, 'h10014c, 'h1001ab, 'h1001ac, 'h1001ae, 'h1001af, 'h100149, 'h10014a, 'h10014b, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b8, 'h10003c, 'h2004f8, 'h100047, 'h1001b7, 'h1001b9, 'h10014c, 'h1001ba, 'h1001bc, 'h1001bb, 'h1001bd, 'h1001be, 'h1001c0, 'h100149, 'h10014a, 'h1001bf, 'h10014b, 'h1001c1, 'h1001c2, 'h1001c4, 'h1001c3, 'h1001c5, 'h10003c, 'h2004f8, 'h100047, 'h1001c6, 'h1001c8, 'h10014c, 'h1001c7, 'h1001c9, 'h1001ca, 'h1001cc, 'h1001cb, 'h1001cd, 'h1001ce, 'h1001d0, 'h1001cf, 'h100149, 'h10014a, 'h10014b, 'h1001d1, 'h1001d3, 'h1001d4, 'h10003c, 'h2004f8, 'h100047, 'h1001d5, 'h1001d7, 'h10014c, 'h1001d8, 'h1001d9, 'h1001db, 'h1001dc, 'h1001dd, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e3, 'h1001e4, 'h100149, 'h10014a, 'h10014b, 'h1001e5, 'h1001e7, 'h1001e8, 'h10003c, 'h2004f8, 'h100047, 'h1001e9, 'h10014c, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f7, 'h1001f8, 'h100149, 'h10014a, 'h10014b, 'h1001f9, 'h1001fb, 'h1001fc, 'h10003c, 'h2004f8, 'h100047, 'h10014c, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h100149, 'h10014a, 'h10014b, 'h10020d, 'h10020f, 'h100210, 'h10003c, 'h2004f8, 'h100047, 'h10014c, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100149, 'h10014a, 'h10014b, 'h100221, 'h100223, 'h100224, 'h10003c, 'h2004f8, 'h100047, 'h10014c, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h100149, 'h10014a, 'h10014b, 'h100235, 'h10003c, 'h2004f8, 'h100047, 'h10014c, 'h100236, 'h100237, 'h100239, 'h100238, 'h10023a, 'h10023b, 'h10023d, 'h10023c, 'h10023e, 'h10023f, 'h100241, 'h100240, 'h100242, 'h100243, 'h100245, 'h100149, 'h10014a, 'h10003c, 'h2004f8, 'h100047, 'h100244, 'h10014b, 'h10014c, 'h100246, 'h100247, 'h100249, 'h100248, 'h10024a, 'h10024b, 'h10024d, 'h10024c, 'h10024e, 'h10024f, 'h100251, 'h100250, 'h100252, 'h100254, 'h100255, 'h10003c, 'h2004f8, 'h100047, 'h100149, 'h10014a, 'h10014b, 'h100256, 'h10014c, 'h100258, 'h100259, 'h10025a, 'h10025c, 'h10025d, 'h10025e, 'h100260, 'h100261, 'h100262, 'h100264, 'h100265, 'h100266, 'h100268, 'h100269, 'h10003c, 'h2004f8, 'h100047, 'h100149, 'h10014a, 'h10014b, 'h10026a, 'h10014c, 'h10026c, 'h10026d, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100150, 'h10014e, 'h100173, 'h10014f, 'h100174, 'h100176, 'h10003c, 'h2004f8, 'h100047, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100186, 'h100150, 'h10014e, 'h100187, 'h10014f, 'h100188, 'h10018a, 'h10003c, 'h2004f8, 'h100047, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h10019a, 'h100150, 'h10014e, 'h10019b, 'h10014f, 'h10019c, 'h10019e, 'h10003c, 'h2004f8, 'h100047, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h100150, 'h10014e, 'h1001af, 'h10014f, 'h1001b0, 'h1001b1, 'h10003c, 'h2004f8, 'h100047, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h100150, 'h1001be, 'h10014e, 'h1001bf, 'h10014f, 'h1001c0, 'h10003c, 'h2004f8, 'h100047, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001ca, 'h1001cb, 'h1001cc, 'h100150, 'h1001cd, 'h1001cf, 'h10014e, 'h1001d0, 'h10014f, 'h10003c, 'h2004f8, 'h100047, 'h1001d1, 'h1001d3, 'h1001d4, 'h1001d5, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001db, 'h1001dc, 'h1001dd, 'h1001df, 'h1001e0, 'h1001e1, 'h100150, 'h1001e3, 'h10014e, 'h1001e4, 'h10014f, 'h10003c, 'h2004f8, 'h100047, 'h1001e5, 'h1001e7, 'h1001e8, 'h1001e9, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h1001f5, 'h100150, 'h1001f7, 'h10014e, 'h1001f8, 'h10014f, 'h10003c, 'h2004f8, 'h100047, 'h1001f9, 'h1001fb, 'h1001fc, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h100150, 'h10020b, 'h10014e, 'h10020c, 'h10014f, 'h10003c, 'h2004f8, 'h100047, 'h10020d, 'h10020f, 'h100210, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h100150, 'h10021f, 'h10014e, 'h100220, 'h10014f, 'h10003c, 'h2004f8, 'h100047, 'h100221, 'h100223, 'h100224, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100150, 'h100232, 'h100233, 'h10014e, 'h100234, 'h10003c, 'h2004f8, 'h100047, 'h10014f, 'h100235, 'h100236, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100150, 'h100242, 'h100243, 'h10014e, 'h10003c, 'h2004f8, 'h100047, 'h100244, 'h10014f, 'h100245, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024b, 'h10024c, 'h10024d, 'h10024e, 'h100250, 'h100251, 'h100252, 'h100150, 'h100254, 'h10014e, 'h10003c, 'h2004f8, 'h100047, 'h100255, 'h10014f, 'h100256, 'h100258, 'h100259, 'h10025a, 'h10025c, 'h10025d, 'h10025e, 'h100260, 'h100261, 'h100262, 'h100264, 'h100265, 'h100266, 'h100150, 'h100268, 'h10014e, 'h10003c, 'h2004f8, 'h100047, 'h100269, 'h10014f, 'h10026a, 'h10026c, 'h10026d, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100154, 'h100152, 'h100173, 'h100153, 'h100174, 'h100176, 'h100177, 'h100178, 'h10003c, 'h2004f8, 'h100047, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100186, 'h100154, 'h100152, 'h100187, 'h100153, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10003c, 'h2004f8, 'h100047, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h10019a, 'h100154, 'h100152, 'h10019b, 'h100153, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h10003c, 'h2004f8, 'h100047, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h100154, 'h100152, 'h1001af, 'h100153, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h10003c, 'h2004f8, 'h100047, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h100154, 'h1001be, 'h100152, 'h1001bf, 'h100153, 'h1001c0, 'h1001c1, 'h1001c2, 'h10003c, 'h2004f8, 'h100047, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c6, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001cb, 'h1001cc, 'h1001cd, 'h100154, 'h1001cf, 'h100152, 'h1001d0, 'h100153, 'h1001d1, 'h1001d3, 'h1001d4, 'h10003c, 'h2004f8, 'h100047, 'h1001d5, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001db, 'h1001dc, 'h1001dd, 'h1001df, 'h1001e0, 'h1001e1, 'h100154, 'h1001e3, 'h100152, 'h1001e4, 'h100153, 'h1001e5, 'h1001e7, 'h1001e8, 'h10003c, 'h2004f8, 'h100047, 'h1001e9, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h1001f5, 'h100154, 'h1001f7, 'h100152, 'h1001f8, 'h100153, 'h1001f9, 'h1001fb, 'h1001fc, 'h10003c, 'h2004f8, 'h100047, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h100154, 'h10020b, 'h100152, 'h10020c, 'h100153, 'h10020d, 'h10020f, 'h100210, 'h10003c, 'h2004f8, 'h100047, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h100154, 'h10021f, 'h100152, 'h100220, 'h100153, 'h100221, 'h100223, 'h100224, 'h10003c, 'h2004f8, 'h100047, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100154, 'h100232, 'h100233, 'h100152, 'h100234, 'h100153, 'h100235, 'h100236, 'h10003c, 'h2004f8, 'h100047, 'h100237, 'h100238, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100154, 'h100242, 'h100243, 'h100152, 'h100244, 'h100153, 'h100245, 'h10003c, 'h2004f8, 'h100047, 'h100246, 'h100247, 'h100248, 'h100249, 'h10024a, 'h10024c, 'h10024d, 'h10024e, 'h100250, 'h100251, 'h100252, 'h100154, 'h100254, 'h100255, 'h100256, 'h100258, 'h100152, 'h100259, 'h10003c, 'h2004f8, 'h100047, 'h100153, 'h10025a, 'h10025c, 'h10025d, 'h10025e, 'h100260, 'h100261, 'h100262, 'h100264, 'h100265, 'h100266, 'h100154, 'h100268, 'h100269, 'h10026a, 'h10026c, 'h100152, 'h10026d, 'h10003c, 'h2004f8, 'h100047, 'h100153, 'h10026e, 'h100270, 'h100271, 'h100272, 'h100172, 'h100158, 'h100156, 'h100173, 'h100157, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10003c, 'h2004f8, 'h100047, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100186, 'h100158, 'h100156, 'h100187, 'h100157, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h10003c, 'h2004f8, 'h100047, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h10019a, 'h100158, 'h100156, 'h10019b, 'h100157, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h10003c, 'h2004f8, 'h100047, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h100158, 'h100156, 'h1001af, 'h100157, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h10003c, 'h2004f8, 'h100047, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h100158, 'h1001be, 'h100156, 'h1001bf, 'h100157, 'h1001c0, 'h1001c1, 'h1001c2, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c7, 'h10003c, 'h2004f8, 'h100047, 'h1001c8, 'h1001c9, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001cf, 'h100158, 'h1001d0, 'h1001d1, 'h1001d3, 'h100156, 'h100157, 'h1001d4, 'h1001d5, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001db, 'h10003c, 'h2004f8, 'h100047, 'h1001dc, 'h1001dd, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e3, 'h100158, 'h1001e4, 'h1001e5, 'h1001e7, 'h100156, 'h1001e8, 'h100157, 'h1001e9, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ef, 'h10003c, 'h2004f8, 'h100047, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f7, 'h100158, 'h1001f8, 'h1001f9, 'h1001fb, 'h100156, 'h1001fc, 'h100157, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h10003c, 'h2004f8, 'h100047, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h100158, 'h10020c, 'h10020d, 'h10020f, 'h100156, 'h100210, 'h100157, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h10003c, 'h2004f8, 'h100047, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100158, 'h100220, 'h100221, 'h100223, 'h100156, 'h100224, 'h100157, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10003c, 'h2004f8, 'h100047, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100158, 'h100233, 'h100234, 'h100235, 'h100236, 'h100237, 'h100156, 'h100238, 'h100157, 'h100239, 'h10023a, 'h10023b, 'h10003c, 'h2004f8, 'h100047, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100158, 'h100242, 'h100243, 'h100244, 'h100245, 'h100246, 'h100248, 'h100156, 'h100157, 'h100249, 'h10024a, 'h10024c, 'h10003c, 'h2004f8, 'h100047, 'h10024d, 'h10024e, 'h100250, 'h100251, 'h100252, 'h100254, 'h100158, 'h100255, 'h100256, 'h100258, 'h100259, 'h10025a, 'h10025c, 'h100156, 'h10025d, 'h100157, 'h10025e, 'h100260, 'h10003c, 'h2004f8, 'h100047, 'h100261, 'h100262, 'h100264, 'h100265, 'h100266, 'h100268, 'h100158, 'h100269, 'h10026a, 'h10026c, 'h10026d, 'h10026e, 'h100270, 'h100156, 'h100271, 'h100157, 'h100272, 'h100172, 'h10015c, 'h10003c, 'h2004f8, 'h100047, 'h10015a, 'h100173, 'h10015b, 'h100174, 'h100176, 'h100177, 'h100178, 'h10017a, 'h10017b, 'h10017c, 'h10017e, 'h10017f, 'h100180, 'h100182, 'h100183, 'h100184, 'h100186, 'h10015c, 'h10003c, 'h2004f8, 'h100047, 'h10015a, 'h100187, 'h10015b, 'h100188, 'h10018a, 'h10018b, 'h10018c, 'h10018e, 'h10018f, 'h100190, 'h100192, 'h100193, 'h100194, 'h100196, 'h100197, 'h100198, 'h10019a, 'h10015c, 'h10003c, 'h2004f8, 'h100047, 'h10015a, 'h10019b, 'h10015b, 'h10019c, 'h10019e, 'h10019f, 'h1001a0, 'h1001a2, 'h1001a3, 'h1001a4, 'h1001a6, 'h1001a7, 'h1001a8, 'h1001aa, 'h1001ab, 'h1001ac, 'h1001ae, 'h10015c, 'h10003c, 'h2004f8, 'h100047, 'h10015a, 'h1001af, 'h10015b, 'h1001b0, 'h1001b1, 'h1001b2, 'h1001b3, 'h1001b4, 'h1001b5, 'h1001b6, 'h1001b7, 'h1001b8, 'h1001b9, 'h1001ba, 'h1001bb, 'h1001bc, 'h1001bd, 'h10015c, 'h10003c, 'h2004f8, 'h100047, 'h1001be, 'h1001bf, 'h10015a, 'h10015b, 'h1001c0, 'h1001c1, 'h1001c3, 'h1001c4, 'h1001c5, 'h1001c7, 'h1001c8, 'h1001c9, 'h1001cb, 'h1001cc, 'h1001cd, 'h1001cf, 'h1001d0, 'h10015c, 'h10003c, 'h2004f8, 'h100047, 'h1001d1, 'h1001d3, 'h10015a, 'h10015b, 'h1001d4, 'h1001d5, 'h1001d7, 'h1001d8, 'h1001d9, 'h1001db, 'h1001dc, 'h1001dd, 'h1001df, 'h1001e0, 'h1001e1, 'h1001e3, 'h1001e4, 'h1001e5, 'h10003c, 'h2004f8, 'h100047, 'h10015c, 'h1001e7, 'h10015a, 'h1001e8, 'h10015b, 'h1001e9, 'h1001eb, 'h1001ec, 'h1001ed, 'h1001ef, 'h1001f0, 'h1001f1, 'h1001f3, 'h1001f4, 'h1001f5, 'h1001f7, 'h1001f8, 'h1001f9, 'h10003c, 'h2004f8, 'h100047, 'h10015c, 'h1001fb, 'h10015a, 'h1001fc, 'h10015b, 'h1001fd, 'h1001ff, 'h100200, 'h100201, 'h100203, 'h100204, 'h100205, 'h100207, 'h100208, 'h100209, 'h10020b, 'h10020c, 'h10020d, 'h10003c, 'h2004f8, 'h100047, 'h10015c, 'h10020f, 'h10015a, 'h100210, 'h10015b, 'h100211, 'h100213, 'h100214, 'h100215, 'h100217, 'h100218, 'h100219, 'h10021b, 'h10021c, 'h10021d, 'h10021f, 'h100220, 'h100221, 'h10003c, 'h2004f8, 'h100047, 'h10015c, 'h100223, 'h10015a, 'h100224, 'h10015b, 'h100225, 'h100227, 'h100228, 'h100229, 'h10022b, 'h10022c, 'h10022d, 'h10022f, 'h100230, 'h100231, 'h100232, 'h100233, 'h100234, 'h10003c, 'h2004f8, 'h100047, 'h100235, 'h10015c, 'h100236, 'h100237, 'h10015a, 'h100238, 'h10015b, 'h100239, 'h10023a, 'h10023b, 'h10023c, 'h10023d, 'h10023e, 'h10023f, 'h100240, 'h100241, 'h100242, 'h100244, 'h10003c, 'h2004f8, 'h100047, 'h100245, 'h10015c, 'h100246, 'h100248, 'h10015a};
	int DATA4 [4*SIZE-1:0] = {DATA3, DATA0};
	
endpackage
