

package LU_PKG;
	
	import LU_PKG_4::DATA4;
	
	parameter LU_DATA_SIZE = 41832, SIZE_LIMIT = 8500;
	
	int DATA0 [LU_DATA_SIZE-(4*SIZE_LIMIT)-1:0] = {'h10249, 'h1015b, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h1003c, 'h204f8, 'h10047, 'h10259, 'h1015c, 'h1025a, 'h1025c, 'h1015a, 'h1025d, 'h1015b, 'h1025e, 'h10260, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1003c, 'h204f8, 'h10047, 'h1026d, 'h1026e, 'h1015c, 'h10270, 'h1015a, 'h10271, 'h1015b, 'h10272, 'h10172, 'h10160, 'h1015e, 'h10173, 'h1015f, 'h10174, 'h10176, 'h10177, 'h10178, 'h1017a, 'h1003c, 'h204f8, 'h10047, 'h1017b, 'h1017c, 'h1017e, 'h1017f, 'h10180, 'h10182, 'h10183, 'h10184, 'h10186, 'h10160, 'h1015e, 'h10187, 'h1015f, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h1003c, 'h204f8, 'h10047, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10196, 'h10197, 'h10198, 'h1019a, 'h10160, 'h1015e, 'h1019b, 'h1015f, 'h1019c, 'h1019e, 'h1019f, 'h101a0, 'h101a2, 'h1003c, 'h204f8, 'h10047, 'h101a3, 'h101a4, 'h101a6, 'h101a7, 'h101a8, 'h101aa, 'h101ab, 'h101ac, 'h101ae, 'h10160, 'h1015e, 'h101af, 'h1015f, 'h101b0, 'h101b1, 'h101b2, 'h101b3, 'h101b4, 'h1003c, 'h204f8, 'h10047, 'h101b5, 'h101b6, 'h101b7, 'h101b8, 'h101b9, 'h101ba, 'h101bb, 'h101bc, 'h101bd, 'h10160, 'h101bf, 'h1015e, 'h1015f, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h101c5, 'h1003c, 'h204f8, 'h10047, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h10160, 'h101d3, 'h1015e, 'h1015f, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h1003c, 'h204f8, 'h10047, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h10160, 'h101e7, 'h1015e, 'h101e8, 'h1015f, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h1003c, 'h204f8, 'h10047, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h10160, 'h101fb, 'h1015e, 'h101fc, 'h1015f, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h1003c, 'h204f8, 'h10047, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h1020d, 'h10160, 'h1020f, 'h1015e, 'h10210, 'h1015f, 'h10211, 'h10213, 'h10214, 'h10215, 'h1003c, 'h204f8, 'h10047, 'h10217, 'h10218, 'h10219, 'h1021b, 'h1021c, 'h1021d, 'h1021f, 'h10220, 'h10221, 'h10160, 'h10223, 'h1015e, 'h10224, 'h1015f, 'h10225, 'h10227, 'h10228, 'h10229, 'h1003c, 'h204f8, 'h10047, 'h1022b, 'h1022c, 'h1022d, 'h1022f, 'h10230, 'h10231, 'h10232, 'h10233, 'h10234, 'h10235, 'h10160, 'h10236, 'h10237, 'h1015e, 'h10238, 'h1015f, 'h10239, 'h1023a, 'h1003c, 'h204f8, 'h10047, 'h1023b, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10160, 'h10248, 'h10249, 'h1024a, 'h1024c, 'h1015e, 'h1015f, 'h1024d, 'h1003c, 'h204f8, 'h10047, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h10160, 'h1025c, 'h1025d, 'h1025e, 'h10260, 'h1015e, 'h10261, 'h1015f, 'h1003c, 'h204f8, 'h10047, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10160, 'h10270, 'h10271, 'h10272, 'h10172, 'h10164, 'h10162, 'h10173, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h10174, 'h10176, 'h10177, 'h10178, 'h1017a, 'h1017b, 'h1017c, 'h1017e, 'h1017f, 'h10180, 'h10182, 'h10183, 'h10184, 'h10186, 'h10164, 'h10162, 'h10187, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10196, 'h10197, 'h10198, 'h1019a, 'h10164, 'h10162, 'h1019b, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h1019c, 'h1019e, 'h1019f, 'h101a0, 'h101a2, 'h101a3, 'h101a4, 'h101a6, 'h101a7, 'h101a8, 'h101aa, 'h101ab, 'h101ac, 'h101ae, 'h10164, 'h10162, 'h101af, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h101b0, 'h101b1, 'h101b2, 'h101b3, 'h101b4, 'h101b5, 'h101b6, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h10164, 'h10162, 'h101c0, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h101c1, 'h101c3, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h10164, 'h10162, 'h101d4, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h10164, 'h10162, 'h101e8, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h10164, 'h10162, 'h101fc, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h1020d, 'h1020f, 'h10164, 'h10162, 'h10210, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h10211, 'h10213, 'h10214, 'h10215, 'h10217, 'h10218, 'h10219, 'h1021b, 'h1021c, 'h1021d, 'h1021f, 'h10220, 'h10221, 'h10223, 'h10164, 'h10162, 'h10224, 'h1003c, 'h204f8, 'h10047, 'h10163, 'h10225, 'h10227, 'h10228, 'h10229, 'h1022b, 'h1022c, 'h1022d, 'h1022f, 'h10230, 'h10231, 'h10232, 'h10233, 'h10234, 'h10235, 'h10164, 'h10236, 'h10237, 'h1003c, 'h204f8, 'h10047, 'h10238, 'h10162, 'h10163, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10164, 'h10249, 'h1024a, 'h1003c, 'h204f8, 'h10047, 'h1024c, 'h10162, 'h10163, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h10164, 'h1025d, 'h1025e, 'h1003c, 'h204f8, 'h10047, 'h10260, 'h10162, 'h10163, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h10164, 'h10271, 'h10272, 'h1003c, 'h204f8, 'h10047, 'h10172, 'h10168, 'h10166, 'h10173, 'h10167, 'h10174, 'h10176, 'h10177, 'h10178, 'h1017a, 'h1017b, 'h1017c, 'h1017e, 'h1017f, 'h10180, 'h10182, 'h10183, 'h10184, 'h1003c, 'h204f8, 'h10047, 'h10186, 'h10168, 'h10166, 'h10187, 'h10167, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10196, 'h10197, 'h10198, 'h1003c, 'h204f8, 'h10047, 'h1019a, 'h10168, 'h10166, 'h1019b, 'h10167, 'h1019c, 'h1019e, 'h1019f, 'h101a0, 'h101a2, 'h101a3, 'h101a4, 'h101a6, 'h101a7, 'h101a8, 'h101aa, 'h101ab, 'h101ac, 'h1003c, 'h204f8, 'h10047, 'h101ae, 'h10168, 'h10166, 'h101af, 'h10167, 'h101b0, 'h101b1, 'h101b2, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h1003c, 'h204f8, 'h10047, 'h101c0, 'h10168, 'h101c1, 'h101c3, 'h10166, 'h10167, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h1003c, 'h204f8, 'h10047, 'h101d4, 'h10168, 'h101d5, 'h101d7, 'h10166, 'h10167, 'h101d8, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h1003c, 'h204f8, 'h10047, 'h101e8, 'h101e9, 'h10168, 'h101eb, 'h10166, 'h101ec, 'h10167, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h1003c, 'h204f8, 'h10047, 'h101fc, 'h101fd, 'h10168, 'h101ff, 'h10166, 'h10200, 'h10167, 'h10201, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h1020d, 'h1020f, 'h1003c, 'h204f8, 'h10047, 'h10210, 'h10211, 'h10168, 'h10213, 'h10166, 'h10214, 'h10167, 'h10215, 'h10217, 'h10218, 'h10219, 'h1021b, 'h1021c, 'h1021d, 'h1021f, 'h10220, 'h10221, 'h10223, 'h1003c, 'h204f8, 'h10047, 'h10224, 'h10225, 'h10168, 'h10227, 'h10166, 'h10228, 'h10167, 'h10229, 'h1022b, 'h1022c, 'h1022d, 'h1022f, 'h10230, 'h10231, 'h10232, 'h10233, 'h10234, 'h10235, 'h1003c, 'h204f8, 'h10047, 'h10236, 'h10238, 'h10168, 'h10239, 'h1023a, 'h1023c, 'h10166, 'h10167, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h1003c, 'h204f8, 'h10047, 'h1024a, 'h1024c, 'h10168, 'h1024d, 'h1024e, 'h10250, 'h10166, 'h10167, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1003c, 'h204f8, 'h10047, 'h1025e, 'h10260, 'h10168, 'h10261, 'h10262, 'h10264, 'h10166, 'h10167, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h1003c, 'h204f8, 'h10047, 'h10272, 'h10172, 'h1016c, 'h1016a, 'h10173, 'h1016b, 'h10174, 'h10176, 'h10177, 'h10178, 'h1017a, 'h1017b, 'h1017c, 'h1017e, 'h1017f, 'h10180, 'h10182, 'h10183, 'h1003c, 'h204f8, 'h10047, 'h10184, 'h10186, 'h1016c, 'h1016a, 'h10187, 'h1016b, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10196, 'h10197, 'h1003c, 'h204f8, 'h10047, 'h10198, 'h1019a, 'h1016c, 'h1016a, 'h1019b, 'h1016b, 'h1019c, 'h1019e, 'h1019f, 'h101a0, 'h101a2, 'h101a3, 'h101a4, 'h101a6, 'h101a7, 'h101a8, 'h101aa, 'h101ab, 'h1003c, 'h204f8, 'h10047, 'h101ac, 'h101ae, 'h1016c, 'h101af, 'h1016a, 'h1016b, 'h101b0, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h1003c, 'h204f8, 'h10047, 'h101c0, 'h101c1, 'h1016c, 'h101c3, 'h1016a, 'h1016b, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h1003c, 'h204f8, 'h10047, 'h101d4, 'h101d5, 'h1016c, 'h101d7, 'h1016a, 'h1016b, 'h101d8, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h1003c, 'h204f8, 'h10047, 'h101e8, 'h101e9, 'h1016c, 'h101eb, 'h1016a, 'h101ec, 'h1016b, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h1003c, 'h204f8, 'h10047, 'h101fc, 'h101fd, 'h1016c, 'h101ff, 'h1016a, 'h10200, 'h1016b, 'h10201, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h1020d, 'h1020f, 'h1003c, 'h204f8, 'h10047, 'h10210, 'h10211, 'h1016c, 'h10213, 'h1016a, 'h10214, 'h1016b, 'h10215, 'h10217, 'h10218, 'h10219, 'h1021b, 'h1021c, 'h1021d, 'h1021f, 'h10220, 'h10221, 'h10223, 'h1003c, 'h204f8, 'h10047, 'h10224, 'h10225, 'h1016c, 'h10227, 'h1016a, 'h10228, 'h1016b, 'h10229, 'h1022b, 'h1022c, 'h1022d, 'h1022f, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h1003c, 'h204f8, 'h10047, 'h10238, 'h10239, 'h1016c, 'h1023a, 'h1023c, 'h1016a, 'h1016b, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h1024a, 'h1003c, 'h204f8, 'h10047, 'h1024c, 'h1024d, 'h1016c, 'h1024e, 'h10250, 'h1016a, 'h1016b, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h1003c, 'h204f8, 'h10047, 'h10260, 'h10261, 'h1016c, 'h10262, 'h10264, 'h1016a, 'h1016b, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10272, 'h1003c, 'h204f8, 'h10047, 'h10172, 'h10170, 'h1016e, 'h10173, 'h1016f, 'h10174, 'h10176, 'h10177, 'h10178, 'h1017a, 'h1017b, 'h1017c, 'h1017e, 'h1017f, 'h10180, 'h10182, 'h10183, 'h10184, 'h1003c, 'h204f8, 'h10047, 'h10186, 'h10170, 'h1016e, 'h10187, 'h1016f, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10196, 'h10197, 'h10198, 'h1003c, 'h204f8, 'h10047, 'h1019a, 'h10170, 'h1016e, 'h1019b, 'h1016f, 'h1019c, 'h1019e, 'h1019f, 'h101a0, 'h101a2, 'h101a3, 'h101a4, 'h101a6, 'h101a7, 'h101a8, 'h101aa, 'h101ab, 'h101ac, 'h1003c, 'h204f8, 'h10047, 'h101af, 'h10170, 'h1016e, 'h101b0, 'h1016f, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h1003c, 'h204f8, 'h10047, 'h101c3, 'h10170, 'h1016e, 'h101c4, 'h1016f, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h1003c, 'h204f8, 'h10047, 'h101d7, 'h10170, 'h1016e, 'h101d8, 'h1016f, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h1003c, 'h204f8, 'h10047, 'h101eb, 'h10170, 'h1016e, 'h101ec, 'h1016f, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h101fc, 'h101fd, 'h1003c, 'h204f8, 'h10047, 'h101ff, 'h10170, 'h1016e, 'h10200, 'h1016f, 'h10201, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h1020d, 'h1020f, 'h10210, 'h10211, 'h1003c, 'h204f8, 'h10047, 'h10213, 'h10170, 'h1016e, 'h10214, 'h1016f, 'h10215, 'h10217, 'h10218, 'h10219, 'h1021b, 'h1021c, 'h1021d, 'h1021f, 'h10220, 'h10221, 'h10223, 'h10224, 'h10225, 'h1003c, 'h204f8, 'h10047, 'h10227, 'h10170, 'h1016e, 'h10228, 'h1016f, 'h10229, 'h1022b, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1003c, 'h204f8, 'h10047, 'h1023c, 'h10170, 'h1016e, 'h1023d, 'h1016f, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h1003c, 'h204f8, 'h10047, 'h10250, 'h10170, 'h1016e, 'h10251, 'h1016f, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h10260, 'h10261, 'h10262, 'h1003c, 'h204f8, 'h10047, 'h10264, 'h10170, 'h1016e, 'h10265, 'h1016f, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10272, 'h204f7, 'h10172, 'h10173, 'h1003c, 'h10174, 'h10047, 'h10176, 'h10178, 'h10177, 'h1017a, 'h1017c, 'h1017b, 'h1017e, 'h10180, 'h1017f, 'h10182, 'h10184, 'h10183, 'h10186, 'h10188, 'h10187, 'h204f7, 'h10172, 'h10173, 'h1003c, 'h10174, 'h10047, 'h1018a, 'h1018c, 'h1018b, 'h1018e, 'h10190, 'h1018f, 'h10192, 'h10194, 'h10193, 'h10196, 'h10198, 'h10197, 'h1019a, 'h1019c, 'h1019b, 'h204f7, 'h10172, 'h10173, 'h1003c, 'h10174, 'h10047, 'h1019e, 'h101a0, 'h1019f, 'h101a2, 'h101a4, 'h101a3, 'h101a6, 'h101a8, 'h101a7, 'h101ab, 'h101ac, 'h101af, 'h101b0, 'h101b1, 'h101b3, 'h204f7, 'h101b4, 'h10172, 'h1003c, 'h10173, 'h10047, 'h10174, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h101c5, 'h101c4, 'h101c7, 'h204f7, 'h101c9, 'h10172, 'h1003c, 'h10173, 'h10047, 'h101c8, 'h10174, 'h101cb, 'h101cd, 'h101cc, 'h101cf, 'h101d1, 'h101d0, 'h101d3, 'h101d5, 'h101d4, 'h101d7, 'h101d9, 'h101d8, 'h101db, 'h204f7, 'h101dd, 'h10172, 'h1003c, 'h10173, 'h10047, 'h101dc, 'h10174, 'h101df, 'h101e1, 'h101e0, 'h101e3, 'h101e5, 'h101e4, 'h101e7, 'h101e9, 'h101e8, 'h101eb, 'h101ed, 'h101ec, 'h101ef, 'h204f7, 'h101f1, 'h10172, 'h1003c, 'h10173, 'h10047, 'h101f0, 'h10174, 'h101f3, 'h101f5, 'h101f4, 'h101f7, 'h101f9, 'h101f8, 'h101fb, 'h101fd, 'h101fc, 'h101ff, 'h10201, 'h10200, 'h10203, 'h204f7, 'h10205, 'h10172, 'h1003c, 'h10204, 'h10047, 'h10173, 'h10174, 'h10207, 'h10209, 'h10208, 'h1020b, 'h1020d, 'h1020c, 'h1020f, 'h10211, 'h10210, 'h10213, 'h10215, 'h10214, 'h10217, 'h204f7, 'h10219, 'h10172, 'h1003c, 'h10218, 'h10047, 'h10173, 'h10174, 'h1021b, 'h1021d, 'h1021c, 'h1021f, 'h10221, 'h10220, 'h10223, 'h10225, 'h10224, 'h10227, 'h10229, 'h10228, 'h1022c, 'h204f7, 'h1022d, 'h10172, 'h1003c, 'h10230, 'h10231, 'h10047, 'h10174, 'h10173, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h204f7, 'h10242, 'h10244, 'h10246, 'h1003c, 'h10172, 'h10047, 'h10245, 'h10173, 'h10174, 'h10248, 'h1024a, 'h10249, 'h1024c, 'h1024e, 'h1024d, 'h10250, 'h10252, 'h10251, 'h10254, 'h10256, 'h204f7, 'h10255, 'h10258, 'h1025a, 'h1003c, 'h10172, 'h10047, 'h10259, 'h10173, 'h10174, 'h1025c, 'h1025e, 'h1025d, 'h10260, 'h10262, 'h10261, 'h10264, 'h10266, 'h10265, 'h10268, 'h1026a, 'h204f7, 'h10269, 'h1026c, 'h1026e, 'h1003c, 'h10172, 'h10047, 'h1026d, 'h10173, 'h10174, 'h10270, 'h10272, 'h10271, 'h1017a, 'h10178, 'h10176, 'h1017b, 'h10177, 'h1017c, 'h1017e, 'h1017f, 'h204f7, 'h10180, 'h10182, 'h10183, 'h1003c, 'h10184, 'h10047, 'h10186, 'h10187, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h10178, 'h10176, 'h1018f, 'h10177, 'h10190, 'h10192, 'h10193, 'h204f7, 'h10194, 'h10196, 'h10197, 'h1003c, 'h10198, 'h10047, 'h1019a, 'h1019b, 'h1019c, 'h1019e, 'h1019f, 'h101a0, 'h101a2, 'h10178, 'h101a3, 'h10176, 'h10177, 'h101a4, 'h101a7, 'h101a8, 'h204f7, 'h101ab, 'h101ac, 'h101af, 'h1003c, 'h101b0, 'h10047, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h10178, 'h101bb, 'h10176, 'h10177, 'h101bc, 'h101bd, 'h101bf, 'h204f7, 'h101c0, 'h101c1, 'h101c3, 'h1003c, 'h101c4, 'h10047, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h10178, 'h101cf, 'h10176, 'h10177, 'h101d0, 'h101d1, 'h101d3, 'h204f7, 'h101d4, 'h101d5, 'h101d7, 'h1003c, 'h101d8, 'h10047, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h10178, 'h101e3, 'h10176, 'h10177, 'h101e4, 'h101e5, 'h101e7, 'h204f7, 'h101e8, 'h101e9, 'h101eb, 'h1003c, 'h101ec, 'h10047, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h10178, 'h101f7, 'h10176, 'h101f8, 'h10177, 'h101f9, 'h101fb, 'h204f7, 'h101fc, 'h101fd, 'h101ff, 'h1003c, 'h10200, 'h10047, 'h10201, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h10178, 'h1020b, 'h10176, 'h1020c, 'h10177, 'h1020d, 'h1020f, 'h204f7, 'h10210, 'h10211, 'h10213, 'h1003c, 'h10214, 'h10047, 'h10215, 'h10217, 'h10218, 'h10219, 'h1021b, 'h1021c, 'h1021d, 'h10178, 'h1021f, 'h10176, 'h10220, 'h10177, 'h10221, 'h10223, 'h204f7, 'h10224, 'h10225, 'h10228, 'h1003c, 'h10229, 'h10047, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10178, 'h10236, 'h10238, 'h10176, 'h10177, 'h10239, 'h1023a, 'h204f7, 'h1023c, 'h1023d, 'h1023e, 'h1003c, 'h10240, 'h10047, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h10178, 'h1024a, 'h1024c, 'h10176, 'h10177, 'h1024d, 'h1024e, 'h204f7, 'h10250, 'h10251, 'h10252, 'h1003c, 'h10254, 'h10047, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h10178, 'h1025e, 'h10260, 'h10176, 'h10177, 'h10261, 'h10262, 'h204f7, 'h10264, 'h10265, 'h10266, 'h1003c, 'h10268, 'h10047, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10178, 'h10272, 'h1017e, 'h1017c, 'h1017a, 'h1017f, 'h1017b, 'h204f7, 'h10180, 'h10182, 'h10183, 'h1003c, 'h10184, 'h10047, 'h10186, 'h10187, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h1017c, 'h1017a, 'h10193, 'h1017b, 'h204f7, 'h10194, 'h10196, 'h10197, 'h1003c, 'h10198, 'h10047, 'h1019a, 'h1019b, 'h1019c, 'h1019e, 'h1019f, 'h101a0, 'h101a3, 'h101a4, 'h101a7, 'h101a8, 'h1017c, 'h101ab, 'h1017a, 'h1017b, 'h204f7, 'h101ac, 'h101af, 'h101b0, 'h1003c, 'h101b1, 'h10047, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h1017c, 'h101c0, 'h101c1, 'h101c3, 'h204f7, 'h1017a, 'h1017b, 'h101c4, 'h1003c, 'h101c5, 'h10047, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h1017c, 'h101d4, 'h101d5, 'h101d7, 'h204f7, 'h1017a, 'h1017b, 'h101d8, 'h1003c, 'h101d9, 'h10047, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h1017c, 'h101e8, 'h101e9, 'h101eb, 'h204f7, 'h1017a, 'h1017b, 'h101ec, 'h1003c, 'h101ed, 'h10047, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h1017c, 'h101fc, 'h101fd, 'h101ff, 'h204f7, 'h1017a, 'h10200, 'h1017b, 'h1003c, 'h10201, 'h10047, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h1020d, 'h1020f, 'h1017c, 'h10210, 'h10211, 'h10213, 'h204f7, 'h1017a, 'h10214, 'h1017b, 'h1003c, 'h10215, 'h10047, 'h10217, 'h10218, 'h10219, 'h1021b, 'h1021c, 'h1021d, 'h1021f, 'h10220, 'h10221, 'h10224, 'h1017c, 'h10225, 'h10228, 'h10229, 'h204f7, 'h1022c, 'h1017a, 'h1017b, 'h1003c, 'h1022d, 'h10047, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1017c, 'h1023d, 'h1023e, 'h10240, 'h204f7, 'h10241, 'h10242, 'h10244, 'h1003c, 'h1017a, 'h10047, 'h1017b, 'h10245, 'h10246, 'h10248, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h1017c, 'h10251, 'h10252, 'h10254, 'h204f7, 'h10255, 'h10256, 'h10258, 'h1003c, 'h1017a, 'h10047, 'h1017b, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h10260, 'h10261, 'h10262, 'h10264, 'h1017c, 'h10265, 'h10266, 'h10268, 'h204f7, 'h10269, 'h1026a, 'h1026c, 'h1003c, 'h1017a, 'h10047, 'h1017b, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10272, 'h10182, 'h10180, 'h1017e, 'h10183, 'h1017f, 'h10184, 'h10186, 'h10187, 'h204f7, 'h10188, 'h1018a, 'h1018b, 'h1003c, 'h1018c, 'h10047, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10196, 'h10180, 'h1017e, 'h10197, 'h1017f, 'h10198, 'h1019a, 'h1019b, 'h204f7, 'h1019c, 'h1019f, 'h101a0, 'h1003c, 'h101a3, 'h10047, 'h101a4, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h101af, 'h101b0, 'h10180, 'h101b1, 'h101b3, 'h1017e, 'h1017f, 'h101b4, 'h101b5, 'h204f7, 'h101b7, 'h101b8, 'h101b9, 'h1003c, 'h101bb, 'h10047, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h10180, 'h101c5, 'h101c7, 'h1017e, 'h1017f, 'h101c8, 'h101c9, 'h204f7, 'h101cb, 'h101cc, 'h101cd, 'h1003c, 'h101cf, 'h10047, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h10180, 'h101d9, 'h101db, 'h1017e, 'h1017f, 'h101dc, 'h101dd, 'h204f7, 'h101df, 'h101e0, 'h101e1, 'h1003c, 'h101e3, 'h10047, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101eb, 'h101ec, 'h10180, 'h101ed, 'h101ef, 'h1017e, 'h1017f, 'h101f0, 'h101f1, 'h204f7, 'h101f3, 'h101f4, 'h101f5, 'h1003c, 'h101f7, 'h10047, 'h101f8, 'h101f9, 'h101fb, 'h101fc, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h10180, 'h10203, 'h1017e, 'h10204, 'h1017f, 'h10205, 'h204f7, 'h10207, 'h10208, 'h10209, 'h1003c, 'h1020b, 'h10047, 'h1020c, 'h1020d, 'h1020f, 'h10210, 'h10211, 'h10213, 'h10214, 'h10215, 'h10180, 'h10217, 'h1017e, 'h10218, 'h1017f, 'h10219, 'h204f7, 'h1021b, 'h1021c, 'h1021d, 'h1003c, 'h10220, 'h10047, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10180, 'h10231, 'h10232, 'h10234, 'h1017e, 'h1017f, 'h204f7, 'h10235, 'h10236, 'h10238, 'h1003c, 'h10239, 'h10047, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10180, 'h10245, 'h10246, 'h10248, 'h1017e, 'h1017f, 'h204f7, 'h10249, 'h1024a, 'h1024c, 'h1003c, 'h1024d, 'h10047, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10180, 'h10259, 'h1025a, 'h1025c, 'h1017e, 'h1017f, 'h204f7, 'h1025d, 'h1025e, 'h10260, 'h1003c, 'h10261, 'h10047, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h10180, 'h1026d, 'h1026e, 'h10270, 'h1017e, 'h1017f, 'h204f7, 'h10271, 'h10272, 'h10186, 'h10184, 'h1003c, 'h10047, 'h10182, 'h10187, 'h10183, 'h10188, 'h1018a, 'h1018b, 'h1018c, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10196, 'h204f7, 'h10197, 'h10198, 'h1019b, 'h10184, 'h1003c, 'h10047, 'h10182, 'h1019c, 'h10183, 'h1019f, 'h101a0, 'h101a3, 'h101a4, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h101af, 'h101b0, 'h101b1, 'h204f7, 'h101b3, 'h101b4, 'h101b5, 'h10184, 'h1003c, 'h10047, 'h101b7, 'h10182, 'h10183, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h101c5, 'h204f7, 'h101c7, 'h101c8, 'h101c9, 'h10184, 'h1003c, 'h10047, 'h101cb, 'h10182, 'h10183, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h204f7, 'h101db, 'h101dc, 'h101dd, 'h10184, 'h1003c, 'h10047, 'h101df, 'h10182, 'h10183, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h204f7, 'h101ef, 'h101f0, 'h101f1, 'h10184, 'h1003c, 'h10047, 'h101f3, 'h10182, 'h10183, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h101fc, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h204f7, 'h10203, 'h10204, 'h10205, 'h10184, 'h1003c, 'h10047, 'h10207, 'h10182, 'h10208, 'h10183, 'h10209, 'h1020b, 'h1020c, 'h1020d, 'h1020f, 'h10210, 'h10211, 'h10213, 'h10214, 'h10215, 'h204f7, 'h10217, 'h10218, 'h10219, 'h10184, 'h1003c, 'h10047, 'h1021c, 'h10182, 'h1021d, 'h10183, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h204f7, 'h10232, 'h10234, 'h10235, 'h10184, 'h1003c, 'h10047, 'h10236, 'h10238, 'h10182, 'h10183, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h204f7, 'h10246, 'h10248, 'h10249, 'h10184, 'h1003c, 'h10047, 'h1024a, 'h1024c, 'h10182, 'h10183, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h204f7, 'h1025a, 'h1025c, 'h1025d, 'h10184, 'h1003c, 'h10047, 'h1025e, 'h10260, 'h10182, 'h10183, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h204f7, 'h1026e, 'h10270, 'h10271, 'h10184, 'h1003c, 'h10047, 'h10272, 'h1018a, 'h10188, 'h10186, 'h1018b, 'h10187, 'h1018c, 'h1018e, 'h1018f, 'h10190, 'h10192, 'h10193, 'h10194, 'h10197, 'h204f7, 'h10198, 'h1019b, 'h1019c, 'h1019f, 'h1003c, 'h10047, 'h101a0, 'h101a3, 'h10188, 'h10186, 'h101a4, 'h10187, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h101af, 'h101b0, 'h101b1, 'h101b3, 'h204f7, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h1003c, 'h10047, 'h101b9, 'h101bb, 'h10188, 'h10186, 'h101bc, 'h10187, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h101c5, 'h101c7, 'h204f7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h1003c, 'h10047, 'h101cd, 'h101cf, 'h10188, 'h10186, 'h101d0, 'h10187, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h101db, 'h204f7, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h1003c, 'h10047, 'h101e1, 'h101e3, 'h10188, 'h10186, 'h101e4, 'h10187, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h101ef, 'h204f7, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h1003c, 'h10047, 'h101f5, 'h101f7, 'h10188, 'h10186, 'h101f8, 'h10187, 'h101f9, 'h101fb, 'h101fc, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h10203, 'h204f7, 'h10204, 'h10205, 'h10207, 'h10208, 'h1003c, 'h10047, 'h10209, 'h1020b, 'h10188, 'h10186, 'h1020c, 'h10187, 'h1020d, 'h1020f, 'h10210, 'h10211, 'h10213, 'h10214, 'h10215, 'h10218, 'h204f7, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h1003c, 'h10047, 'h10221, 'h10224, 'h10188, 'h10186, 'h10225, 'h10187, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h204f7, 'h10235, 'h10236, 'h10238, 'h10239, 'h1003c, 'h10047, 'h1023a, 'h1023c, 'h10188, 'h10186, 'h1023d, 'h10187, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h204f7, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1003c, 'h10047, 'h1024e, 'h10250, 'h10188, 'h10186, 'h10251, 'h10187, 'h10252, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h204f7, 'h1025d, 'h1025e, 'h10260, 'h10261, 'h1003c, 'h10047, 'h10262, 'h10264, 'h10188, 'h10186, 'h10265, 'h10187, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h204f7, 'h10271, 'h10272, 'h1018e, 'h1018c, 'h1018f, 'h1003c, 'h10047, 'h1018a, 'h1018b, 'h10190, 'h10193, 'h10194, 'h10197, 'h10198, 'h1019b, 'h1019c, 'h1019f, 'h101a0, 'h101a3, 'h101a4, 'h204f7, 'h101a7, 'h101a8, 'h101ab, 'h1018c, 'h101ac, 'h1003c, 'h10047, 'h101af, 'h1018a, 'h1018b, 'h101b0, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h204f7, 'h101bd, 'h101bf, 'h101c0, 'h1018c, 'h101c1, 'h1003c, 'h10047, 'h101c3, 'h1018a, 'h1018b, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h204f7, 'h101d1, 'h101d3, 'h101d4, 'h1018c, 'h101d5, 'h1003c, 'h10047, 'h101d7, 'h1018a, 'h1018b, 'h101d8, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h204f7, 'h101e5, 'h101e7, 'h101e8, 'h1018c, 'h101e9, 'h1003c, 'h10047, 'h101eb, 'h101ec, 'h1018a, 'h1018b, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h204f7, 'h101f9, 'h101fb, 'h101fc, 'h1018c, 'h101fd, 'h1003c, 'h10047, 'h101ff, 'h10200, 'h1018a, 'h1018b, 'h10201, 'h10203, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h204f7, 'h1020d, 'h1020f, 'h10210, 'h1018c, 'h10211, 'h1003c, 'h10047, 'h10214, 'h10215, 'h10218, 'h1018a, 'h1018b, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h204f7, 'h10229, 'h1022c, 'h1022d, 'h1018c, 'h10230, 'h1003c, 'h10047, 'h10231, 'h10232, 'h10234, 'h1018a, 'h1018b, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h204f7, 'h10240, 'h10241, 'h10242, 'h1018c, 'h10244, 'h1003c, 'h10047, 'h10245, 'h10246, 'h10248, 'h1018a, 'h1018b, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h204f7, 'h10254, 'h10255, 'h10256, 'h1018c, 'h10258, 'h1003c, 'h10047, 'h10259, 'h1025a, 'h1025c, 'h1018a, 'h1018b, 'h1025d, 'h1025e, 'h10260, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h204f7, 'h10268, 'h10269, 'h1026a, 'h1018c, 'h1026c, 'h1026d, 'h1003c, 'h10047, 'h1026e, 'h10270, 'h10271, 'h1018a, 'h1018b, 'h10272, 'h10193, 'h10190, 'h1018f, 'h10194, 'h10197, 'h10198, 'h204f7, 'h1019b, 'h1019c, 'h1019f, 'h101a0, 'h101a3, 'h101a4, 'h1003c, 'h10047, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h101af, 'h101b0, 'h101b1, 'h10190, 'h101b3, 'h1018f, 'h101b4, 'h101b5, 'h204f7, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h1003c, 'h10047, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h101c5, 'h101c7, 'h10190, 'h101c8, 'h1018f, 'h101c9, 'h101cb, 'h204f7, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h1003c, 'h10047, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h101db, 'h101dc, 'h10190, 'h101dd, 'h101df, 'h1018f, 'h101e0, 'h204f7, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h1003c, 'h10047, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h10190, 'h101f3, 'h101f4, 'h1018f, 'h101f5, 'h204f7, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h101fc, 'h101fd, 'h1003c, 'h10047, 'h101ff, 'h10200, 'h10201, 'h10203, 'h10204, 'h10205, 'h10207, 'h10190, 'h10208, 'h10209, 'h1020b, 'h1020c, 'h1018f, 'h204f7, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h1003c, 'h10047, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10190, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1018f, 'h204f7, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h1003c, 'h10047, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h10190, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h204f7, 'h1018f, 'h10245, 'h10246, 'h10248, 'h10249, 'h1003c, 'h10047, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10190, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h204f7, 'h1018f, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h1003c, 'h10047, 'h10260, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10190, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h204f7, 'h10270, 'h1018f, 'h10271, 'h10272, 'h10197, 'h10194, 'h1003c, 'h10047, 'h10193, 'h10198, 'h1019b, 'h1019c, 'h1019f, 'h101a0, 'h101a3, 'h101a4, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h204f7, 'h101af, 'h101b0, 'h101b1, 'h101b3, 'h101b4, 'h10194, 'h1003c, 'h10047, 'h101b5, 'h101b7, 'h10193, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h204f7, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h10194, 'h1003c, 'h10047, 'h101cb, 'h101cc, 'h10193, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h204f7, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h10194, 'h1003c, 'h10047, 'h101e0, 'h101e1, 'h101e3, 'h10193, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h204f7, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h10194, 'h1003c, 'h10047, 'h101f5, 'h101f7, 'h101f8, 'h10193, 'h101f9, 'h101fb, 'h101fc, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h10203, 'h204f7, 'h10204, 'h10205, 'h10207, 'h10208, 'h10209, 'h10194, 'h1003c, 'h10047, 'h1020c, 'h1020d, 'h10210, 'h10193, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h204f7, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h10194, 'h1003c, 'h10047, 'h1022c, 'h1022d, 'h10230, 'h10193, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h204f7, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10194, 'h1003c, 'h10047, 'h10242, 'h10244, 'h10245, 'h10193, 'h10246, 'h10248, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h204f7, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h10194, 'h1003c, 'h10047, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h10193, 'h1025d, 'h1025e, 'h10260, 'h10261, 'h10262, 'h10264, 'h10265, 'h204f7, 'h10266, 'h10268, 'h10269, 'h1026a, 'h1026c, 'h10194, 'h1003c, 'h10047, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10193, 'h10272, 'h1019b, 'h10198, 'h10197, 'h1019c, 'h1019f, 'h101a0, 'h204f7, 'h101a3, 'h101a4, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h1003c, 'h10047, 'h101af, 'h101b0, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h10198, 'h10197, 'h101b8, 'h101b9, 'h101bb, 'h204f7, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h1003c, 'h10047, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h10198, 'h101cd, 'h101cf, 'h10197, 'h101d0, 'h204f7, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h1003c, 'h10047, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h10198, 'h101e3, 'h101e4, 'h10197, 'h101e5, 'h204f7, 'h101e7, 'h101e8, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h1003c, 'h10047, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h10198, 'h101f8, 'h101f9, 'h101fb, 'h101fc, 'h204f7, 'h10197, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h10203, 'h10204, 'h1003c, 'h10047, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10198, 'h10211, 'h10214, 'h10215, 'h10218, 'h204f7, 'h10197, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h1003c, 'h10047, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10198, 'h10231, 'h10232, 'h10234, 'h10235, 'h204f7, 'h10197, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1003c, 'h10047, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10198, 'h10246, 'h10248, 'h10249, 'h1024a, 'h204f7, 'h1024c, 'h10197, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h1003c, 'h10047, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h10198, 'h1025c, 'h1025d, 'h1025e, 'h10260, 'h204f7, 'h10261, 'h10197, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1003c, 'h10047, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h10198, 'h10271, 'h10272, 'h1019f, 'h1019c, 'h204f7, 'h1019b, 'h101a0, 'h101a3, 'h101a4, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h1003c, 'h10047, 'h101af, 'h101b0, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h1019c, 'h204f7, 'h101bb, 'h1019b, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h1003c, 'h10047, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h1019c, 'h204f7, 'h101d0, 'h1019b, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h1003c, 'h10047, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h1019c, 'h204f7, 'h101e5, 'h101e7, 'h1019b, 'h101e8, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h1003c, 'h10047, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h1019c, 'h204f7, 'h101fb, 'h101fc, 'h1019b, 'h101fd, 'h101ff, 'h10200, 'h10201, 'h10204, 'h1003c, 'h10047, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h1019c, 'h204f7, 'h10218, 'h10219, 'h1021c, 'h1019b, 'h1021d, 'h10220, 'h10221, 'h10224, 'h1003c, 'h10047, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h1019c, 'h204f7, 'h10235, 'h10236, 'h10238, 'h1019b, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1003c, 'h10047, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h1019c, 'h204f7, 'h1024a, 'h1024c, 'h1024d, 'h1019b, 'h1024e, 'h10250, 'h10251, 'h10252, 'h1003c, 'h10047, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h1019c, 'h204f7, 'h10260, 'h10261, 'h10262, 'h10264, 'h1019b, 'h10265, 'h10266, 'h10268, 'h1003c, 'h10047, 'h10269, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10272, 'h101a3, 'h101a0, 'h204f7, 'h1019f, 'h101a4, 'h101a7, 'h101a8, 'h101ab, 'h101ac, 'h101af, 'h101b0, 'h1003c, 'h10047, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101a0, 'h204f7, 'h101bd, 'h101bf, 'h1019f, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h101c5, 'h1003c, 'h10047, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101a0, 'h204f7, 'h101d3, 'h101d4, 'h1019f, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h101db, 'h1003c, 'h10047, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101a0, 'h204f7, 'h101e8, 'h101e9, 'h101eb, 'h1019f, 'h101ec, 'h101ed, 'h101ef, 'h101f0, 'h1003c, 'h10047, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h101f8, 'h101f9, 'h101fb, 'h101fc, 'h101a0, 'h204f7, 'h101fd, 'h10200, 'h10201, 'h10204, 'h1019f, 'h10205, 'h10208, 'h10209, 'h1003c, 'h10047, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h101a0, 'h204f7, 'h1021d, 'h10220, 'h10221, 'h10224, 'h1019f, 'h10225, 'h10228, 'h10229, 'h1003c, 'h10047, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h101a0, 'h204f7, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1019f, 'h1023e, 'h10240, 'h10241, 'h1003c, 'h10047, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h101a0, 'h204f7, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h1019f, 'h10255, 'h10256, 'h1003c, 'h10047, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h10260, 'h10261, 'h10262, 'h101a0, 'h204f7, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1019f, 'h1026a, 'h1026c, 'h1003c, 'h10047, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10272, 'h101a7, 'h101a4, 'h101a3, 'h101a8, 'h101ab, 'h204f7, 'h101ac, 'h101af, 'h101b0, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h1003c, 'h10047, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101a4, 'h101a3, 'h101c0, 'h101c1, 'h204f7, 'h101c3, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h1003c, 'h10047, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101a4, 'h101d5, 'h101d7, 'h101a3, 'h204f7, 'h101d8, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h1003c, 'h10047, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101a4, 'h101eb, 'h101ec, 'h101a3, 'h204f7, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h101f7, 'h1003c, 'h10047, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h101a4, 'h10204, 'h10205, 'h10208, 'h204f7, 'h101a3, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h1003c, 'h10047, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h101a4, 'h10224, 'h10225, 'h10228, 'h204f7, 'h101a3, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h1003c, 'h10047, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h101a4, 'h1023d, 'h1023e, 'h10240, 'h204f7, 'h101a3, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h1003c, 'h10047, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h101a4, 'h10252, 'h10254, 'h10255, 'h204f7, 'h101a3, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h1003c, 'h10047, 'h10260, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h101a4, 'h10268, 'h10269, 'h1026a, 'h204f7, 'h1026c, 'h101a3, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10272, 'h101ab, 'h101a8, 'h1003c, 'h10047, 'h101a7, 'h101ac, 'h101ad, 'h101af, 'h101b0, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h204f7, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101a8, 'h1003c, 'h10047, 'h101c1, 'h101c3, 'h101a7, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h204f7, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101a8, 'h1003c, 'h10047, 'h101d7, 'h101d8, 'h101a7, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h204f7, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101eb, 'h101a8, 'h1003c, 'h10047, 'h101ec, 'h101ed, 'h101ef, 'h101a7, 'h101f0, 'h101f1, 'h101f3, 'h101f4, 'h101f5, 'h204f7, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h101a8, 'h1003c, 'h10047, 'h10208, 'h10209, 'h1020c, 'h101a7, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h204f7, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h101a8, 'h1003c, 'h10047, 'h10228, 'h10229, 'h1022c, 'h101a7, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h204f7, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h101a8, 'h1003c, 'h10047, 'h10240, 'h10241, 'h10242, 'h10244, 'h101a7, 'h10245, 'h10246, 'h10248, 'h10249, 'h204f7, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h101a8, 'h1003c, 'h10047, 'h10255, 'h10256, 'h10258, 'h10259, 'h101a7, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h204f7, 'h10260, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h101a8, 'h1003c, 'h10047, 'h1026a, 'h1026c, 'h1026d, 'h1026e, 'h10270, 'h101a7, 'h10271, 'h10272, 'h101af, 'h204f7, 'h101ad, 'h101ab, 'h101b0, 'h101ac, 'h101b1, 'h101b3, 'h101b4, 'h101b5, 'h101b7, 'h1003c, 'h10047, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h204f7, 'h101ad, 'h101ab, 'h101c4, 'h101ac, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h1003c, 'h10047, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h204f7, 'h101ad, 'h101ab, 'h101d8, 'h101ac, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h1003c, 'h10047, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101eb, 'h204f7, 'h101ad, 'h101ab, 'h101ec, 'h101ac, 'h101ed, 'h101ef, 'h101f0, 'h101f1, 'h101f4, 'h1003c, 'h10047, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h204f7, 'h10208, 'h101ad, 'h101ab, 'h101ac, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h1003c, 'h10047, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h204f7, 'h10225, 'h10228, 'h101ad, 'h101ab, 'h101ac, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h1003c, 'h10047, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h204f7, 'h1023d, 'h1023e, 'h10240, 'h101ad, 'h101ab, 'h10241, 'h101ac, 'h10242, 'h10244, 'h1003c, 'h10047, 'h10245, 'h10246, 'h10248, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h204f7, 'h10251, 'h10252, 'h10254, 'h101ad, 'h101ab, 'h10255, 'h101ac, 'h10256, 'h10258, 'h1003c, 'h10047, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h10260, 'h10261, 'h10262, 'h10264, 'h204f7, 'h10265, 'h10266, 'h10268, 'h101ad, 'h101ab, 'h10269, 'h101ac, 'h1026a, 'h1026c, 'h1003c, 'h10047, 'h1026d, 'h1026e, 'h10270, 'h10271, 'h10272, 'h101b3, 'h101b1, 'h101af, 'h101b4, 'h204f7, 'h101b0, 'h101b5, 'h101b7, 'h101b8, 'h101b9, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h1003c, 'h10047, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h101c5, 'h101c7, 'h101b1, 'h101af, 'h101c8, 'h204f7, 'h101b0, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h1003c, 'h10047, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h101db, 'h101b1, 'h101dc, 'h101af, 'h204f7, 'h101b0, 'h101dd, 'h101df, 'h101e0, 'h101e1, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h1003c, 'h10047, 'h101e9, 'h101eb, 'h101ec, 'h101ed, 'h101f0, 'h101b1, 'h101f1, 'h101f4, 'h204f7, 'h101af, 'h101b0, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h1003c, 'h10047, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h101b1, 'h10210, 'h10211, 'h204f7, 'h10214, 'h101af, 'h101b0, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h1003c, 'h10047, 'h10224, 'h10225, 'h10228, 'h10229, 'h1022c, 'h101b1, 'h1022d, 'h10230, 'h204f7, 'h10231, 'h10232, 'h10234, 'h101af, 'h10235, 'h101b0, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1003c, 'h10047, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h101b1, 'h10244, 'h204f7, 'h10245, 'h10246, 'h10248, 'h101af, 'h10249, 'h101b0, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h1003c, 'h10047, 'h10250, 'h10251, 'h10252, 'h10254, 'h10255, 'h10256, 'h101b1, 'h10258, 'h204f7, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h101af, 'h101b0, 'h1025e, 'h10260, 'h10261, 'h10262, 'h1003c, 'h10047, 'h10264, 'h10265, 'h10266, 'h10268, 'h10269, 'h1026a, 'h101b1, 'h1026c, 'h204f7, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h101b7, 'h101b5, 'h101b3, 'h101b8, 'h101b4, 'h101b9, 'h1003c, 'h10047, 'h101bb, 'h101bc, 'h101bd, 'h101bf, 'h101c0, 'h101c1, 'h101c3, 'h101c4, 'h204f7, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101b5, 'h101b3, 'h101cc, 'h101b4, 'h101cd, 'h1003c, 'h10047, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h204f7, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101b5, 'h101b3, 'h101e0, 'h101b4, 'h101e1, 'h1003c, 'h10047, 'h101e3, 'h101e4, 'h101e5, 'h101e7, 'h101e8, 'h101e9, 'h101ec, 'h101ed, 'h204f7, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101b5, 'h101b3, 'h101f9, 'h101b4, 'h101fc, 'h1003c, 'h10047, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h1020c, 'h204f7, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h101b5, 'h10218, 'h101b3, 'h101b4, 'h10219, 'h1003c, 'h10047, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h204f7, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h101b5, 'h10234, 'h101b3, 'h10235, 'h101b4, 'h1003c, 'h10047, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h204f7, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h101b5, 'h10248, 'h101b3, 'h10249, 'h101b4, 'h1003c, 'h10047, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h10254, 'h204f7, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h101b5, 'h1025c, 'h101b3, 'h1025d, 'h101b4, 'h1003c, 'h10047, 'h1025e, 'h10260, 'h10261, 'h10262, 'h10264, 'h10265, 'h10266, 'h10268, 'h204f7, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h101b5, 'h10272, 'h101bb, 'h101b9, 'h101bd, 'h1003c, 'h10047, 'h101b7, 'h101bc, 'h101b8, 'h101bf, 'h101c1, 'h101c0, 'h101c3, 'h101c5, 'h204f7, 'h101c4, 'h101c7, 'h101c9, 'h101c8, 'h101cb, 'h101cd, 'h101cc, 'h101cf, 'h101b9, 'h101d1, 'h1003c, 'h10047, 'h101b7, 'h101d0, 'h101b8, 'h101d3, 'h101d5, 'h101d4, 'h101d7, 'h101d9, 'h204f7, 'h101d8, 'h101db, 'h101dd, 'h101dc, 'h101df, 'h101e1, 'h101e0, 'h101e3, 'h101b9, 'h101e5, 'h1003c, 'h10047, 'h101e4, 'h101b7, 'h101b8, 'h101e8, 'h101e9, 'h101ec, 'h101ed, 'h101f0, 'h204f7, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h101b9, 'h10201, 'h1003c, 'h10047, 'h10204, 'h10205, 'h101b7, 'h101b8, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h204f7, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h101b9, 'h10220, 'h10221, 'h1003c, 'h10047, 'h10224, 'h10225, 'h101b7, 'h101b8, 'h10228, 'h10229, 'h1022c, 'h204f7, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10236, 'h10235, 'h10238, 'h101b9, 'h1023a, 'h10239, 'h1003c, 'h10047, 'h1023c, 'h1023e, 'h101b7, 'h1023d, 'h101b8, 'h10240, 'h10242, 'h204f7, 'h10241, 'h10244, 'h10246, 'h10245, 'h10248, 'h1024a, 'h10249, 'h1024c, 'h101b9, 'h1024e, 'h1024d, 'h1003c, 'h10047, 'h10250, 'h10252, 'h101b7, 'h10251, 'h101b8, 'h10254, 'h10256, 'h204f7, 'h10255, 'h10258, 'h1025a, 'h10259, 'h1025c, 'h1025e, 'h1025d, 'h10260, 'h101b9, 'h10262, 'h10261, 'h1003c, 'h10047, 'h10264, 'h10266, 'h10265, 'h101b7, 'h101b8, 'h10269, 'h1026a, 'h204f7, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h101bf, 'h101bd, 'h101bb, 'h101c0, 'h101bc, 'h101c1, 'h101c3, 'h1003c, 'h10047, 'h101c4, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h204f7, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101bd, 'h101bb, 'h101d4, 'h101bc, 'h101d5, 'h101d7, 'h1003c, 'h10047, 'h101d8, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101df, 'h101e0, 'h204f7, 'h101e1, 'h101e4, 'h101e5, 'h101e8, 'h101e9, 'h101bd, 'h101ec, 'h101bb, 'h101bc, 'h101ed, 'h101f0, 'h1003c, 'h10047, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h204f7, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h101bd, 'h10209, 'h1020c, 'h101bb, 'h101bc, 'h1020d, 'h1003c, 'h10047, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h204f7, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h101bd, 'h10228, 'h10229, 'h1022c, 'h101bb, 'h101bc, 'h1003c, 'h10047, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h204f7, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h101bd, 'h10240, 'h10241, 'h101bb, 'h101bc, 'h1003c, 'h10047, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h10249, 'h1024a, 'h204f7, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h101bd, 'h10254, 'h10255, 'h101bb, 'h101bc, 'h1003c, 'h10047, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h204f7, 'h10260, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h101bd, 'h1026a, 'h1026d, 'h101bb, 'h101bc, 'h1003c, 'h10047, 'h1026e, 'h10271, 'h10272, 'h101c3, 'h101c1, 'h101c4, 'h101bf, 'h204f7, 'h101c0, 'h101c5, 'h101c7, 'h101c8, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h1003c, 'h10047, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101c1, 'h101d8, 'h101bf, 'h204f7, 'h101c0, 'h101d9, 'h101db, 'h101dc, 'h101dd, 'h101e0, 'h101e1, 'h101e4, 'h101e5, 'h101e8, 'h101e9, 'h1003c, 'h10047, 'h101ec, 'h101ed, 'h101f0, 'h101f1, 'h101c1, 'h101f4, 'h101bf, 'h204f7, 'h101c0, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h1003c, 'h10047, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h101c1, 'h10211, 'h10214, 'h204f7, 'h101bf, 'h101c0, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h1003c, 'h10047, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h101c1, 'h10230, 'h10231, 'h204f7, 'h101bf, 'h101c0, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1003c, 'h10047, 'h1023e, 'h10240, 'h10241, 'h10242, 'h101c1, 'h10244, 'h10245, 'h204f7, 'h101bf, 'h101c0, 'h10246, 'h10248, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h1003c, 'h10047, 'h10252, 'h10254, 'h10255, 'h10256, 'h101c1, 'h10258, 'h10259, 'h204f7, 'h101bf, 'h101c0, 'h1025a, 'h1025c, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1003c, 'h10047, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h101c1, 'h10272, 'h101c7, 'h204f7, 'h101c5, 'h101c3, 'h101c8, 'h101c4, 'h101c9, 'h101cb, 'h101cc, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h1003c, 'h10047, 'h101d3, 'h101d4, 'h101d5, 'h101d7, 'h101d8, 'h101d9, 'h101dc, 'h204f7, 'h101c5, 'h101c3, 'h101dd, 'h101c4, 'h101e0, 'h101e1, 'h101e4, 'h101e5, 'h101e8, 'h101e9, 'h101ec, 'h1003c, 'h10047, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h204f7, 'h101c5, 'h101fc, 'h101c3, 'h101c4, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h1003c, 'h10047, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h204f7, 'h101c5, 'h10219, 'h1021c, 'h101c3, 'h101c4, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h1003c, 'h10047, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h204f7, 'h101c5, 'h10235, 'h10236, 'h10238, 'h101c3, 'h101c4, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h1003c, 'h10047, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h204f7, 'h101c5, 'h10249, 'h1024a, 'h1024c, 'h101c3, 'h1024d, 'h101c4, 'h1024e, 'h10250, 'h10251, 'h10252, 'h1003c, 'h10047, 'h10254, 'h10255, 'h10256, 'h10258, 'h10259, 'h1025a, 'h1025d, 'h204f7, 'h101c5, 'h1025e, 'h10261, 'h10262, 'h10265, 'h101c3, 'h101c4, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1003c, 'h10047, 'h1026e, 'h10271, 'h10272, 'h101cb, 'h101c9, 'h101c7, 'h101cc, 'h204f7, 'h101c8, 'h101cd, 'h101cf, 'h101d0, 'h101d1, 'h101d3, 'h101d4, 'h101d5, 'h101d8, 'h101d9, 'h101dc, 'h1003c, 'h10047, 'h101dd, 'h101e0, 'h101e1, 'h101e4, 'h101c9, 'h101c7, 'h101e5, 'h204f7, 'h101c8, 'h101e8, 'h101e9, 'h101ec, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h1003c, 'h10047, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h101c9, 'h10204, 'h101c7, 'h204f7, 'h101c8, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h1003c, 'h10047, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h101c9, 'h10221, 'h10224, 'h204f7, 'h101c7, 'h101c8, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h1003c, 'h10047, 'h10235, 'h10236, 'h10238, 'h10239, 'h101c9, 'h1023a, 'h1023c, 'h204f7, 'h101c7, 'h101c8, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h1003c, 'h10047, 'h10249, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h101c9, 'h10250, 'h204f7, 'h101c7, 'h10251, 'h101c8, 'h10252, 'h10254, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h1003c, 'h10047, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h101c9, 'h1026a, 'h204f7, 'h1026d, 'h101c7, 'h101c8, 'h1026e, 'h10271, 'h10272, 'h101cf, 'h101cd, 'h101d0, 'h101cb, 'h101cc, 'h1003c, 'h10047, 'h101d1, 'h101d4, 'h101d5, 'h101d8, 'h101d9, 'h101dc, 'h101dd, 'h204f7, 'h101e0, 'h101e1, 'h101e4, 'h101e5, 'h101e8, 'h101e9, 'h101ec, 'h101cd, 'h101ed, 'h101f0, 'h101cb, 'h1003c, 'h10047, 'h101cc, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h204f7, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h101cd, 'h1020c, 'h1020d, 'h10210, 'h1003c, 'h10047, 'h101cb, 'h101cc, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h204f7, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h101cd, 'h10229, 'h1022c, 'h1022d, 'h1003c, 'h10047, 'h10230, 'h101cb, 'h101cc, 'h10231, 'h10232, 'h10234, 'h10235, 'h204f7, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h101cd, 'h10240, 'h10241, 'h10242, 'h1003c, 'h10047, 'h10244, 'h10245, 'h101cb, 'h101cc, 'h10246, 'h10248, 'h10249, 'h204f7, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10250, 'h10251, 'h10252, 'h101cd, 'h10255, 'h10256, 'h10259, 'h1003c, 'h10047, 'h1025a, 'h1025d, 'h101cb, 'h101cc, 'h1025e, 'h10261, 'h10262, 'h204f7, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h101cd, 'h10272, 'h101d4, 'h101d1, 'h1003c, 'h10047, 'h101d0, 'h101d5, 'h101d8, 'h101d9, 'h101dc, 'h101dd, 'h101e0, 'h204f7, 'h101e1, 'h101e4, 'h101e5, 'h101e8, 'h101e9, 'h101ec, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h101d1, 'h1003c, 'h10047, 'h101d0, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h204f7, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h101d1, 'h1003c, 'h10047, 'h101d0, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h204f7, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h101d1, 'h1003c, 'h10047, 'h10234, 'h101d0, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h204f7, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h101d1, 'h1003c, 'h10047, 'h10249, 'h101d0, 'h1024a, 'h1024c, 'h1024d, 'h1024e, 'h10251, 'h204f7, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h101d1, 'h1003c, 'h10047, 'h10266, 'h101d0, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h204f7, 'h10272, 'h101d8, 'h101d5, 'h101d9, 'h101d4, 'h101dc, 'h101dd, 'h101e0, 'h101e1, 'h101e4, 'h101e5, 'h1003c, 'h10047, 'h101e8, 'h101e9, 'h101ec, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h204f7, 'h101f5, 'h101f8, 'h101d5, 'h101f9, 'h101d4, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h1003c, 'h10047, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h204f7, 'h10215, 'h10218, 'h101d5, 'h10219, 'h101d4, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h1003c, 'h10047, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h204f7, 'h10234, 'h10235, 'h101d5, 'h10236, 'h10238, 'h10239, 'h101d4, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h1003c, 'h10047, 'h10240, 'h10241, 'h10242, 'h10244, 'h10245, 'h10246, 'h10248, 'h204f7, 'h10249, 'h1024a, 'h101d5, 'h1024d, 'h1024e, 'h10251, 'h101d4, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1003c, 'h10047, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h204f7, 'h10269, 'h1026a, 'h101d5, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h101d4, 'h101dc, 'h101d9, 'h101d8, 'h101dd, 'h1003c, 'h10047, 'h101e0, 'h101e1, 'h101e4, 'h101e5, 'h101e8, 'h101e9, 'h204f7, 'h101ec, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101d9, 'h101d8, 'h101fd, 'h1003c, 'h10047, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h204f7, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h101d9, 'h101d8, 'h1021d, 'h1003c, 'h10047, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h204f7, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h101d9, 'h101d8, 'h10239, 'h1003c, 'h10047, 'h1023a, 'h1023c, 'h1023d, 'h1023e, 'h10240, 'h10241, 'h204f7, 'h10242, 'h10244, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h101d9, 'h101d8, 'h10252, 'h1003c, 'h10047, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h204f7, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h101d9, 'h101d8, 'h10272, 'h1003c, 'h10047, 'h101e0, 'h101dd, 'h101dc, 'h101e1, 'h101e4, 'h101e5, 'h204f7, 'h101e8, 'h101e9, 'h101ec, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h1003c, 'h10047, 'h10200, 'h101dd, 'h101dc, 'h10201, 'h10204, 'h10205, 'h204f7, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h1003c, 'h10047, 'h10220, 'h101dd, 'h101dc, 'h10221, 'h10224, 'h10225, 'h204f7, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1003c, 'h10047, 'h1023a, 'h101dd, 'h1023c, 'h1023d, 'h101dc, 'h1023e, 'h204f7, 'h10240, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h1003c, 'h10047, 'h10256, 'h101dd, 'h10259, 'h1025a, 'h1025d, 'h101dc, 'h204f7, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h101e4, 'h101e1, 'h1003c, 'h10047, 'h101e0, 'h101e5, 'h101e8, 'h101e9, 'h101ec, 'h204f7, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h101e1, 'h1003c, 'h10047, 'h101e0, 'h10205, 'h10208, 'h10209, 'h1020c, 'h204f7, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h101e1, 'h1003c, 'h10047, 'h101e0, 'h10225, 'h10228, 'h10229, 'h1022c, 'h204f7, 'h1022d, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023c, 'h1023d, 'h101e1, 'h1003c, 'h10047, 'h1023e, 'h10241, 'h101e0, 'h10242, 'h10245, 'h204f7, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h101e1, 'h1003c, 'h10047, 'h1025e, 'h10261, 'h101e0, 'h10262, 'h10265, 'h204f7, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h101e8, 'h101e5, 'h101e4, 'h101e9, 'h101ec, 'h101ed, 'h1003c, 'h10047, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h204f7, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h101e5, 'h101e4, 'h10209, 'h1020c, 'h1020d, 'h1003c, 'h10047, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h204f7, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h101e5, 'h101e4, 'h10229, 'h1022c, 'h1022d, 'h1003c, 'h10047, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h204f7, 'h10236, 'h10238, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h101e5, 'h10245, 'h101e4, 'h10246, 'h10249, 'h1003c, 'h10047, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h204f7, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h101e5, 'h10265, 'h101e4, 'h10266, 'h10269, 'h1003c, 'h10047, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h204f7, 'h101ec, 'h101e9, 'h101e8, 'h101ed, 'h101f0, 'h101f1, 'h101f4, 'h101f5, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h1003c, 'h10047, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h204f7, 'h1020c, 'h101e9, 'h101e8, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h1003c, 'h10047, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h204f7, 'h1022c, 'h101e9, 'h1022d, 'h101e8, 'h10230, 'h10231, 'h10232, 'h10234, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1003c, 'h10047, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h204f7, 'h10249, 'h101e9, 'h1024a, 'h1024d, 'h101e8, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1003c, 'h10047, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h204f7, 'h10269, 'h101e9, 'h1026a, 'h1026d, 'h101e8, 'h1026e, 'h10271, 'h10272, 'h101f0, 'h101ed, 'h101f1, 'h101ec, 'h101f4, 'h101f5, 'h1003c, 'h10047, 'h101f8, 'h101f9, 'h101fc, 'h101fd, 'h204f7, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h101ed, 'h10211, 'h101ec, 'h10214, 'h10215, 'h1003c, 'h10047, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h204f7, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10230, 'h101ed, 'h10231, 'h101ec, 'h10232, 'h10235, 'h1003c, 'h10047, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h204f7, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h101ed, 'h10251, 'h101ec, 'h10252, 'h10255, 'h1003c, 'h10047, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h204f7, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h101ed, 'h10271, 'h10272, 'h101ec, 'h101f4, 'h101f1, 'h1003c, 'h10047, 'h101f0, 'h101f5, 'h101f8, 'h204f7, 'h101f9, 'h101fc, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h101f1, 'h1003c, 'h10047, 'h101f0, 'h10215, 'h10218, 'h204f7, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h1022c, 'h1022d, 'h10231, 'h10232, 'h10235, 'h101f1, 'h1003c, 'h10047, 'h101f0, 'h10236, 'h10239, 'h204f7, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h101f1, 'h1003c, 'h10047, 'h101f0, 'h10256, 'h10259, 'h204f7, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h101f8, 'h101f5, 'h1003c, 'h10047, 'h101f4, 'h101f9, 'h101fc, 'h204f7, 'h101fd, 'h10200, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h101f5, 'h1003c, 'h10047, 'h101f4, 'h10219, 'h1021c, 'h204f7, 'h1021d, 'h10220, 'h10221, 'h10224, 'h10225, 'h10228, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h101f5, 'h1003c, 'h10047, 'h1023d, 'h101f4, 'h1023e, 'h204f7, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h101f5, 'h1003c, 'h10047, 'h1025d, 'h101f4, 'h1025e, 'h204f7, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h101fc, 'h101f9, 'h101fd, 'h101f8, 'h10200, 'h10201, 'h1003c, 'h10047, 'h10204, 'h10205, 'h204f7, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h101f9, 'h1021d, 'h101f8, 'h10220, 'h10221, 'h1003c, 'h10047, 'h10224, 'h10225, 'h204f7, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h101f9, 'h10242, 'h10245, 'h101f8, 'h10246, 'h1003c, 'h10047, 'h10249, 'h1024a, 'h204f7, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h101f9, 'h10262, 'h10265, 'h10266, 'h101f8, 'h1003c, 'h10047, 'h10269, 'h1026a, 'h204f7, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h10200, 'h101fd, 'h101fc, 'h10201, 'h10204, 'h10205, 'h10208, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h1003c, 'h10047, 'h10214, 'h10215, 'h204f7, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10220, 'h101fd, 'h10221, 'h101fc, 'h10225, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1003c, 'h10047, 'h1023a, 'h1023d, 'h204f7, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h101fd, 'h10249, 'h101fc, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1003c, 'h10047, 'h1025a, 'h1025d, 'h204f7, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h101fd, 'h10269, 'h101fc, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h10204, 'h10201, 'h10205, 'h1003c, 'h10047, 'h10200, 'h10208, 'h204f7, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021c, 'h1021d, 'h10221, 'h10225, 'h10229, 'h10201, 'h1022d, 'h1003c, 'h10047, 'h10200, 'h10231, 'h204f7, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h10201, 'h1024e, 'h1003c, 'h10047, 'h10251, 'h10200, 'h204f7, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h10201, 'h1026e, 'h1003c, 'h10047, 'h10271, 'h10272, 'h204f7, 'h10200, 'h10208, 'h10205, 'h10204, 'h10209, 'h1020c, 'h1020d, 'h10210, 'h10211, 'h10214, 'h10215, 'h10218, 'h10219, 'h1021d, 'h10221, 'h10225, 'h1003c, 'h10047, 'h10229, 'h1022d, 'h204f7, 'h10231, 'h10232, 'h10205, 'h10235, 'h10204, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1003c, 'h10047, 'h1024d, 'h1024e, 'h204f7, 'h10251, 'h10252, 'h10205, 'h10255, 'h10204, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1003c, 'h10047, 'h1026d, 'h1026e, 'h204f7, 'h10271, 'h10272, 'h10205, 'h1020c, 'h10209, 'h1020d, 'h10208, 'h10210, 'h10211, 'h10214, 'h10215, 'h10219, 'h1021d, 'h10221, 'h10225, 'h10229, 'h1003c, 'h10047, 'h1022d, 'h10231, 'h204f7, 'h10232, 'h10235, 'h10236, 'h10239, 'h10209, 'h1023a, 'h1023d, 'h10208, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h1003c, 'h10047, 'h10251, 'h204f7, 'h10252, 'h10255, 'h10256, 'h10259, 'h10209, 'h1025a, 'h1025d, 'h1025e, 'h10208, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h1003c, 'h10047, 'h10271, 'h204f7, 'h10272, 'h10210, 'h1020d, 'h10211, 'h1020c, 'h10215, 'h10219, 'h1021d, 'h10221, 'h10225, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1003c, 'h10047, 'h1023a, 'h204f7, 'h1023d, 'h1023e, 'h1020d, 'h10241, 'h1020c, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1003c, 'h10047, 'h204f7, 'h1025d, 'h1025e, 'h1020d, 'h10261, 'h10262, 'h1020c, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h10215, 'h10211, 'h10219, 'h1021d, 'h1003c, 'h10047, 'h204f7, 'h10221, 'h10225, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10211, 'h10246, 'h10249, 'h1003c, 'h10047, 'h204f7, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10211, 'h10269, 'h1026a, 'h1003c, 'h10047, 'h204f7, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h10219, 'h10215, 'h1021d, 'h10221, 'h10225, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1003c, 'h10047, 'h204f7, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10215, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h1003c, 'h10047, 'h204f7, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h10215, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h1021d, 'h10219, 'h10221, 'h10225, 'h10229, 'h1022d, 'h10231, 'h1003c, 'h10047, 'h204f7, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h10219, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h1003c, 'h10047, 'h204f7, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h10219, 'h1026d, 'h1026e, 'h10271, 'h10272, 'h10221, 'h1021d, 'h1003c, 'h204f7, 'h10047, 'h10225, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1021d, 'h1003c, 'h204f7, 'h10047, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1021d, 'h1003c, 'h204f7, 'h10047, 'h1026e, 'h10271, 'h10272, 'h10225, 'h10221, 'h10229, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h1003c, 'h204f7, 'h10047, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h10221, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h1003c, 'h204f7, 'h10047, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10221, 'h10271, 'h10272, 'h10229, 'h10225, 'h1022d, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h1003c, 'h204f7, 'h10047, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10225, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h1003c, 'h204f7, 'h10047, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10225, 'h10272, 'h1022d, 'h10229, 'h1022e, 'h10231, 'h10232, 'h10235, 'h10236, 'h10239, 'h1003c, 'h204f7, 'h10047, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10229, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1003c, 'h204f7, 'h10047, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h10229, 'h10272, 'h10231, 'h1022e, 'h1022d, 'h10232, 'h10235, 'h1003c, 'h204f7, 'h10047, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h1022e, 'h1022d, 'h10252, 'h10255, 'h1003c, 'h204f7, 'h10047, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10271, 'h1022e, 'h10272, 'h1022d, 'h10235, 'h10232, 'h1003c, 'h204f7, 'h10047, 'h10231, 'h10236, 'h10239, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10232, 'h1003c, 'h204f7, 'h10047, 'h10231, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026d, 'h1026e, 'h10272, 'h10239, 'h10236, 'h10235, 'h1003c, 'h204f7, 'h10047, 'h1023a, 'h1023d, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h10236, 'h10235, 'h1003c, 'h204f7, 'h10047, 'h1025a, 'h1025d, 'h1025e, 'h10261, 'h10262, 'h10265, 'h10266, 'h10269, 'h1026a, 'h1026e, 'h10272, 'h1023d, 'h1023a, 'h10239, 'h1023e, 'h10241, 'h10242, 'h10245, 'h10246, 'h1003c, 'h204f7, 'h10047, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1023a, 'h1025e, 'h10239, 'h10261, 'h10262, 'h10265, 'h10266, 'h1003c, 'h204f7, 'h10047, 'h1026a, 'h1026e, 'h10272, 'h10241, 'h1023e, 'h10242, 'h1023d, 'h10245, 'h10246, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1003c, 'h204f7, 'h10047, 'h1025d, 'h1025e, 'h10261, 'h1023e, 'h10262, 'h1023d, 'h10266, 'h1026a, 'h1026e, 'h10272, 'h10245, 'h10242, 'h10246, 'h10241, 'h10249, 'h1024a, 'h1024d, 'h1024e, 'h1003c, 'h204f7, 'h10047, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025d, 'h1025e, 'h10262, 'h10266, 'h1026a, 'h10242, 'h1026e, 'h10241, 'h10272, 'h10249, 'h10246, 'h10245, 'h1003c, 'h204f7, 'h10047, 'h1024a, 'h1024d, 'h1024e, 'h10251, 'h10252, 'h10255, 'h10256, 'h10259, 'h1025a, 'h1025e, 'h10262, 'h10266, 'h1026a, 'h1026e, 'h10272, 'h10249, 'h204f8, 'h10044, 'h1003e, 'h204f7, 'h1003f, 'h10040, 'h10041, 'h10042, 'h10043};
	int LU_DATA [LU_DATA_SIZE-1:0] = {DATA4, DATA0};
	
endpackage
