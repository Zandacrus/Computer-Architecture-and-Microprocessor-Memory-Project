

package MATRIX_MULTIPLY_16_PKG;
	
	parameter MM16_DATA_SIZE = 9075;
	
	int MM16_DATA [MM16_DATA_SIZE-1:0] = {'h21f91, 'h103be, 'h106b8, 'h21f90, 'h21f8f, 'h21f8d, 'h103c0, 'h21f8a, 'h21f8c, 'h103c1, 'h11f9c, 'h103bc, 'h10005, 'h11f9d, 'h10002, 'h21f8e, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106de, 'h106df, 'h106e0, 'h21f8c, 'h106e1, 'h106e2, 'h103bc, 'h106e3, 'h106e4, 'h106e5, 'h106e6, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h106e7, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106e8, 'h106e9, 'h21f8c, 'h106ea, 'h106eb, 'h103bc, 'h106ec, 'h106ed, 'h106ee, 'h106ef, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h106f0, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106f1, 'h106f2, 'h21f8c, 'h106f3, 'h106f4, 'h103bc, 'h106f5, 'h106f6, 'h106f7, 'h106f8, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h106f9, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h106fa, 'h106fb, 'h21f8c, 'h106fc, 'h106fd, 'h103bc, 'h106fe, 'h106ff, 'h10700, 'h10701, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10702, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10703, 'h10704, 'h21f8c, 'h10705, 'h10706, 'h103bc, 'h10707, 'h10708, 'h10709, 'h1070a, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1070b, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1070c, 'h1070d, 'h21f8c, 'h1070e, 'h1070f, 'h103bc, 'h10710, 'h10711, 'h10712, 'h10713, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10714, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10715, 'h10716, 'h21f8c, 'h10717, 'h10718, 'h103bc, 'h10719, 'h1071a, 'h1071b, 'h1071c, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1071d, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1071e, 'h1071f, 'h21f8c, 'h10720, 'h10721, 'h103bc, 'h10722, 'h10723, 'h10724, 'h10725, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10726, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10727, 'h10728, 'h21f8c, 'h10729, 'h1072a, 'h103bc, 'h1072b, 'h1072c, 'h1072d, 'h1072e, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1072f, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10730, 'h10731, 'h21f8c, 'h10732, 'h10733, 'h103bc, 'h10734, 'h10735, 'h10736, 'h10737, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10738, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10739, 'h1073a, 'h21f8c, 'h1073b, 'h1073c, 'h103bc, 'h1073d, 'h1073e, 'h1073f, 'h10740, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10741, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10742, 'h10743, 'h21f8c, 'h10744, 'h10745, 'h103bc, 'h10746, 'h10747, 'h10748, 'h10749, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1074a, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1074b, 'h1074c, 'h21f8c, 'h1074d, 'h1074e, 'h103bc, 'h1074f, 'h10750, 'h10751, 'h10752, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10753, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10754, 'h10755, 'h21f8c, 'h10756, 'h10757, 'h103bc, 'h10758, 'h10759, 'h1075a, 'h1075b, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1075c, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1075d, 'h21f8d, 'h21f8c, 'h1075e, 'h1075f, 'h103bc, 'h10760, 'h10761, 'h10762, 'h10763, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10764, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10765, 'h10766, 'h21f8c, 'h10767, 'h10768, 'h103bc, 'h10769, 'h1076a, 'h1076b, 'h1076c, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1076d, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1076e, 'h1076f, 'h21f8c, 'h10770, 'h10771, 'h103bc, 'h10772, 'h10773, 'h10774, 'h10775, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10776, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10777, 'h10778, 'h21f8c, 'h10779, 'h1077a, 'h103bc, 'h1077b, 'h1077c, 'h1077d, 'h1077e, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1077f, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10780, 'h10781, 'h21f8c, 'h10782, 'h10783, 'h103bc, 'h10784, 'h10785, 'h10786, 'h10787, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10788, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10789, 'h1078a, 'h21f8c, 'h1078b, 'h1078c, 'h103bc, 'h1078d, 'h1078e, 'h1078f, 'h10790, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h10791, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h10792, 'h10793, 'h21f8c, 'h10794, 'h10795, 'h103bc, 'h10796, 'h10797, 'h10798, 'h10799, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h1079a, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h1079b, 'h1079c, 'h21f8c, 'h1079d, 'h1079e, 'h103bc, 'h1079f, 'h107a0, 'h107a1, 'h107a2, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107a3, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107a4, 'h107a5, 'h21f8c, 'h107a6, 'h107a7, 'h103bc, 'h107a8, 'h107a9, 'h107aa, 'h107ab, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107ac, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107ad, 'h107ae, 'h21f8c, 'h107af, 'h107b0, 'h103bc, 'h107b1, 'h107b2, 'h107b3, 'h107b4, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107b5, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107b6, 'h107b7, 'h21f8c, 'h107b8, 'h107b9, 'h103bc, 'h107ba, 'h107bb, 'h107bc, 'h107bd, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107be, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107bf, 'h107c0, 'h21f8c, 'h107c1, 'h107c2, 'h103bc, 'h107c3, 'h107c4, 'h107c5, 'h107c6, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107c7, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107c8, 'h107c9, 'h21f8c, 'h107ca, 'h107cb, 'h103bc, 'h107cc, 'h107cd, 'h107ce, 'h107cf, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107d0, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107d1, 'h107d2, 'h21f8c, 'h107d3, 'h107d4, 'h103bc, 'h107d5, 'h107d6, 'h107d7, 'h107d8, 'h10001, 'h10000, 'h103bf, 'h21f8b, 'h107d9, 'h21f89, 'h21f83, 'h21f87, 'h21f84, 'h21f85, 'h103b9, 'h107da, 'h107db, 'h21f8c, 'h107dc, 'h107dd, 'h103bc, 'h21f8d, 'h107de, 'h107df, 'h107e0, 'h107e1, 'h107e2, 'h107e3, 'h21f8b, 'h107e4, 'h107e5, 'h107e6, 'h107e7, 'h107e8, 'h107e9, 'h107ea, 'h107eb, 'h107ec, 'h107ed, 'h107ee, 'h107ef, 'h103bc, 'h107f0, 'h107f1, 'h107f2, 'h107f3, 'h107f4, 'h107f5, 'h107f6, 'h21f8b, 'h107f7, 'h107f8, 'h107f9, 'h107fa, 'h107fb, 'h107fc, 'h107fd, 'h107fe, 'h107ff, 'h10800, 'h10801, 'h10802, 'h103bc, 'h10803, 'h10804, 'h10805, 'h10806, 'h10807, 'h10808, 'h10809, 'h21f8b, 'h1080a, 'h1080b, 'h1080c, 'h1080d, 'h1080e, 'h1080f, 'h10810, 'h10811, 'h10812, 'h10813, 'h10814, 'h10815, 'h103bc, 'h10816, 'h10817, 'h10818, 'h10819, 'h1081a, 'h1081b, 'h1081c, 'h21f8b, 'h1081d, 'h1081e, 'h1081f, 'h10820, 'h10821, 'h10822, 'h10823, 'h10824, 'h10825, 'h10826, 'h10827, 'h10828, 'h103bc, 'h10829, 'h1082a, 'h1082b, 'h1082c, 'h1082d, 'h1082e, 'h1082f, 'h21f8b, 'h10830, 'h10831, 'h10832, 'h10833, 'h10834, 'h10835, 'h10836, 'h10837, 'h10838, 'h10839, 'h1083a, 'h1083b, 'h103bc, 'h1083c, 'h1083d, 'h1083e, 'h1083f, 'h10840, 'h10841, 'h10842, 'h21f8b, 'h10843, 'h10844, 'h10845, 'h10846, 'h10847, 'h10848, 'h10849, 'h1084a, 'h1084b, 'h1084c, 'h1084d, 'h1084e, 'h103bc, 'h1084f, 'h10850, 'h10851, 'h10852, 'h10853, 'h10854, 'h10855, 'h21f8b, 'h10856, 'h10857, 'h10858, 'h10859, 'h1085a, 'h1085b, 'h1085c, 'h1085d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1075e, 'h107de, 'h103bc, 'h106e6, 'h106ee, 'h1075f, 'h106f6, 'h106fe, 'h10760, 'h10706, 'h1070e, 'h10761, 'h10716, 'h1071e, 'h10762, 'h10726, 'h1072e, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h107de, 'h103bc, 'h1073e, 'h10764, 'h10746, 'h1074e, 'h10765, 'h10756, 'h106de, 'h10766, 'h107e6, 'h106e6, 'h106ee, 'h10767, 'h106f6, 'h106fe, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10769, 'h103bc, 'h10716, 'h1071e, 'h1076a, 'h10726, 'h1072e, 'h1076b, 'h10736, 'h107e6, 'h1073e, 'h1076c, 'h10746, 'h1074e, 'h1076d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1076e, 'h107ee, 'h103bc, 'h106e6, 'h106ee, 'h1076f, 'h106f6, 'h106fe, 'h10770, 'h10706, 'h1070e, 'h10771, 'h10716, 'h1071e, 'h10772, 'h10726, 'h1072e, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h107ee, 'h103bc, 'h1073e, 'h10774, 'h10746, 'h1074e, 'h10775, 'h10756, 'h106de, 'h10776, 'h107f6, 'h106e6, 'h106ee, 'h10777, 'h106f6, 'h106fe, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10779, 'h103bc, 'h10716, 'h1071e, 'h1077a, 'h10726, 'h1072e, 'h1077b, 'h10736, 'h107f6, 'h1073e, 'h1077c, 'h10746, 'h1074e, 'h1077d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1077e, 'h107fe, 'h103bc, 'h106e6, 'h106ee, 'h1077f, 'h106f6, 'h106fe, 'h10780, 'h10706, 'h1070e, 'h10781, 'h10716, 'h1071e, 'h10782, 'h10726, 'h1072e, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h107fe, 'h103bc, 'h1073e, 'h10784, 'h10746, 'h1074e, 'h10785, 'h10756, 'h106de, 'h10786, 'h10806, 'h106e6, 'h106ee, 'h10787, 'h106f6, 'h106fe, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10789, 'h103bc, 'h10716, 'h1071e, 'h1078a, 'h10726, 'h1072e, 'h1078b, 'h10736, 'h10806, 'h1073e, 'h1078c, 'h10746, 'h1074e, 'h1078d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1078e, 'h1080e, 'h103bc, 'h106e6, 'h106ee, 'h1078f, 'h106f6, 'h106fe, 'h10790, 'h10706, 'h1070e, 'h10791, 'h10716, 'h1071e, 'h10792, 'h10726, 'h1072e, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1080e, 'h103bc, 'h1073e, 'h10794, 'h10746, 'h1074e, 'h10795, 'h10756, 'h106de, 'h10796, 'h10816, 'h106e6, 'h106ee, 'h10797, 'h106f6, 'h106fe, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10799, 'h103bc, 'h10716, 'h1071e, 'h1079a, 'h10726, 'h1072e, 'h1079b, 'h10736, 'h10816, 'h1073e, 'h1079c, 'h10746, 'h1074e, 'h1079d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1079e, 'h1081e, 'h103bc, 'h106e6, 'h106ee, 'h1079f, 'h106f6, 'h106fe, 'h107a0, 'h10706, 'h1070e, 'h107a1, 'h10716, 'h1071e, 'h107a2, 'h10726, 'h1072e, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1081e, 'h103bc, 'h1073e, 'h107a4, 'h10746, 'h1074e, 'h107a5, 'h10756, 'h106de, 'h107a6, 'h10826, 'h106e6, 'h106ee, 'h107a7, 'h106f6, 'h106fe, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107a9, 'h103bc, 'h10716, 'h1071e, 'h107aa, 'h10726, 'h1072e, 'h107ab, 'h10736, 'h10826, 'h1073e, 'h107ac, 'h10746, 'h1074e, 'h107ad, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h107ae, 'h1082e, 'h103bc, 'h106e6, 'h106ee, 'h107af, 'h106f6, 'h106fe, 'h107b0, 'h10706, 'h1070e, 'h107b1, 'h10716, 'h1071e, 'h107b2, 'h10726, 'h1072e, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1082e, 'h103bc, 'h1073e, 'h107b4, 'h10746, 'h1074e, 'h107b5, 'h10756, 'h106de, 'h107b6, 'h10836, 'h106e6, 'h106ee, 'h107b7, 'h106f6, 'h106fe, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107b9, 'h103bc, 'h10716, 'h1071e, 'h107ba, 'h10726, 'h1072e, 'h107bb, 'h10736, 'h10836, 'h1073e, 'h107bc, 'h10746, 'h1074e, 'h107bd, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h107be, 'h1083e, 'h103bc, 'h106e6, 'h106ee, 'h107bf, 'h106f6, 'h106fe, 'h107c0, 'h10706, 'h1070e, 'h107c1, 'h10716, 'h1071e, 'h107c2, 'h10726, 'h1072e, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1083e, 'h103bc, 'h1073e, 'h107c4, 'h10746, 'h1074e, 'h107c5, 'h10756, 'h106de, 'h107c6, 'h10846, 'h106e6, 'h106ee, 'h107c7, 'h106f6, 'h106fe, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107c9, 'h103bc, 'h10716, 'h1071e, 'h107ca, 'h10726, 'h1072e, 'h107cb, 'h10736, 'h10846, 'h1073e, 'h107cc, 'h10746, 'h1074e, 'h107cd, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h107ce, 'h1084e, 'h103bc, 'h106e6, 'h106ee, 'h107cf, 'h106f6, 'h106fe, 'h107d0, 'h10706, 'h1070e, 'h107d1, 'h10716, 'h1071e, 'h107d2, 'h10726, 'h1072e, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1084e, 'h103bc, 'h1073e, 'h107d4, 'h10746, 'h1074e, 'h107d5, 'h10756, 'h106de, 'h107d6, 'h10856, 'h106e6, 'h106ee, 'h107d7, 'h106f6, 'h106fe, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107d9, 'h103bc, 'h10716, 'h1071e, 'h107da, 'h10726, 'h1072e, 'h107db, 'h10736, 'h10856, 'h1073e, 'h107dc, 'h10746, 'h1074e, 'h107dd, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1075e, 'h107de, 'h103bc, 'h106e6, 'h106ee, 'h1075f, 'h106f6, 'h106fe, 'h10760, 'h10706, 'h1070e, 'h10761, 'h10716, 'h1071e, 'h10762, 'h10726, 'h1072e, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h107de, 'h103bc, 'h1073e, 'h10764, 'h10746, 'h1074e, 'h10765, 'h10756, 'h106de, 'h10766, 'h107e6, 'h106e6, 'h106ee, 'h10767, 'h106f6, 'h106fe, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10769, 'h103bc, 'h10716, 'h1071e, 'h1076a, 'h10726, 'h1072e, 'h1076b, 'h10736, 'h107e6, 'h1073e, 'h1076c, 'h10746, 'h1074e, 'h1076d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1076e, 'h107ee, 'h103bc, 'h106e6, 'h106ee, 'h1076f, 'h106f6, 'h106fe, 'h10770, 'h10706, 'h1070e, 'h10771, 'h10716, 'h1071e, 'h10772, 'h10726, 'h1072e, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h107ee, 'h103bc, 'h1073e, 'h10774, 'h10746, 'h1074e, 'h10775, 'h10756, 'h106de, 'h10776, 'h107f6, 'h106e6, 'h106ee, 'h10777, 'h106f6, 'h106fe, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10779, 'h103bc, 'h10716, 'h1071e, 'h1077a, 'h10726, 'h1072e, 'h1077b, 'h10736, 'h107f6, 'h1073e, 'h1077c, 'h10746, 'h1074e, 'h1077d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1077e, 'h107fe, 'h103bc, 'h106e6, 'h106ee, 'h1077f, 'h106f6, 'h106fe, 'h10780, 'h10706, 'h1070e, 'h10781, 'h10716, 'h1071e, 'h10782, 'h10726, 'h1072e, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h107fe, 'h103bc, 'h1073e, 'h10784, 'h10746, 'h1074e, 'h10785, 'h10756, 'h106de, 'h10786, 'h10806, 'h106e6, 'h106ee, 'h10787, 'h106f6, 'h106fe, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10789, 'h103bc, 'h10716, 'h1071e, 'h1078a, 'h10726, 'h1072e, 'h1078b, 'h10736, 'h10806, 'h1073e, 'h1078c, 'h10746, 'h1074e, 'h1078d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1078e, 'h1080e, 'h103bc, 'h106e6, 'h106ee, 'h1078f, 'h106f6, 'h106fe, 'h10790, 'h10706, 'h1070e, 'h10791, 'h10716, 'h1071e, 'h10792, 'h10726, 'h1072e, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1080e, 'h103bc, 'h1073e, 'h10794, 'h10746, 'h1074e, 'h10795, 'h10756, 'h106de, 'h10796, 'h10816, 'h106e6, 'h106ee, 'h10797, 'h106f6, 'h106fe, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h10799, 'h103bc, 'h10716, 'h1071e, 'h1079a, 'h10726, 'h1072e, 'h1079b, 'h10736, 'h10816, 'h1073e, 'h1079c, 'h10746, 'h1074e, 'h1079d, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h1079e, 'h1081e, 'h103bc, 'h106e6, 'h106ee, 'h1079f, 'h106f6, 'h106fe, 'h107a0, 'h10706, 'h1070e, 'h107a1, 'h10716, 'h1071e, 'h107a2, 'h10726, 'h1072e, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1081e, 'h103bc, 'h1073e, 'h107a4, 'h10746, 'h1074e, 'h107a5, 'h10756, 'h106de, 'h107a6, 'h10826, 'h106e6, 'h106ee, 'h107a7, 'h106f6, 'h106fe, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107a9, 'h103bc, 'h10716, 'h1071e, 'h107aa, 'h10726, 'h1072e, 'h107ab, 'h10736, 'h10826, 'h1073e, 'h107ac, 'h10746, 'h1074e, 'h107ad, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h107ae, 'h1082e, 'h103bc, 'h106e6, 'h106ee, 'h107af, 'h106f6, 'h106fe, 'h107b0, 'h10706, 'h1070e, 'h107b1, 'h10716, 'h1071e, 'h107b2, 'h10726, 'h1072e, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1082e, 'h103bc, 'h1073e, 'h107b4, 'h10746, 'h1074e, 'h107b5, 'h10756, 'h106de, 'h107b6, 'h10836, 'h106e6, 'h106ee, 'h107b7, 'h106f6, 'h106fe, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107b9, 'h103bc, 'h10716, 'h1071e, 'h107ba, 'h10726, 'h1072e, 'h107bb, 'h10736, 'h10836, 'h1073e, 'h107bc, 'h10746, 'h1074e, 'h107bd, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h107be, 'h1083e, 'h103bc, 'h106e6, 'h106ee, 'h107bf, 'h106f6, 'h106fe, 'h107c0, 'h10706, 'h1070e, 'h107c1, 'h10716, 'h1071e, 'h107c2, 'h10726, 'h1072e, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1083e, 'h103bc, 'h1073e, 'h107c4, 'h10746, 'h1074e, 'h107c5, 'h10756, 'h106de, 'h107c6, 'h10846, 'h106e6, 'h106ee, 'h107c7, 'h106f6, 'h106fe, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107c9, 'h103bc, 'h10716, 'h1071e, 'h107ca, 'h10726, 'h1072e, 'h107cb, 'h10736, 'h10846, 'h1073e, 'h107cc, 'h10746, 'h1074e, 'h107cd, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106de, 'h107ce, 'h1084e, 'h103bc, 'h106e6, 'h106ee, 'h107cf, 'h106f6, 'h106fe, 'h107d0, 'h10706, 'h1070e, 'h107d1, 'h10716, 'h1071e, 'h107d2, 'h10726, 'h1072e, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h1084e, 'h103bc, 'h1073e, 'h107d4, 'h10746, 'h1074e, 'h107d5, 'h10756, 'h106de, 'h107d6, 'h10856, 'h106e6, 'h106ee, 'h107d7, 'h106f6, 'h106fe, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1070e, 'h107d9, 'h103bc, 'h10716, 'h1071e, 'h107da, 'h10726, 'h1072e, 'h107db, 'h10736, 'h10856, 'h1073e, 'h107dc, 'h10746, 'h1074e, 'h107dd, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1075e, 'h107df, 'h103bc, 'h106e7, 'h106ef, 'h1075f, 'h106f7, 'h106ff, 'h10760, 'h10707, 'h1070f, 'h10761, 'h10717, 'h1071f, 'h10762, 'h10727, 'h1072f, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h107df, 'h103bc, 'h1073f, 'h10764, 'h10747, 'h1074f, 'h10765, 'h10757, 'h106df, 'h10766, 'h107e7, 'h106e7, 'h106ef, 'h10767, 'h106f7, 'h106ff, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10769, 'h103bc, 'h10717, 'h1071f, 'h1076a, 'h10727, 'h1072f, 'h1076b, 'h10737, 'h107e7, 'h1073f, 'h1076c, 'h10747, 'h1074f, 'h1076d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1076e, 'h107ef, 'h103bc, 'h106e7, 'h106ef, 'h1076f, 'h106f7, 'h106ff, 'h10770, 'h10707, 'h1070f, 'h10771, 'h10717, 'h1071f, 'h10772, 'h10727, 'h1072f, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h107ef, 'h103bc, 'h1073f, 'h10774, 'h10747, 'h1074f, 'h10775, 'h10757, 'h106df, 'h10776, 'h107f7, 'h106e7, 'h106ef, 'h10777, 'h106f7, 'h106ff, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10779, 'h103bc, 'h10717, 'h1071f, 'h1077a, 'h10727, 'h1072f, 'h1077b, 'h10737, 'h107f7, 'h1073f, 'h1077c, 'h10747, 'h1074f, 'h1077d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1077e, 'h107ff, 'h103bc, 'h106e7, 'h106ef, 'h1077f, 'h106f7, 'h106ff, 'h10780, 'h10707, 'h1070f, 'h10781, 'h10717, 'h1071f, 'h10782, 'h10727, 'h1072f, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h107ff, 'h103bc, 'h1073f, 'h10784, 'h10747, 'h1074f, 'h10785, 'h10757, 'h106df, 'h10786, 'h10807, 'h106e7, 'h106ef, 'h10787, 'h106f7, 'h106ff, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10789, 'h103bc, 'h10717, 'h1071f, 'h1078a, 'h10727, 'h1072f, 'h1078b, 'h10737, 'h10807, 'h1073f, 'h1078c, 'h10747, 'h1074f, 'h1078d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1078e, 'h1080f, 'h103bc, 'h106e7, 'h106ef, 'h1078f, 'h106f7, 'h106ff, 'h10790, 'h10707, 'h1070f, 'h10791, 'h10717, 'h1071f, 'h10792, 'h10727, 'h1072f, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1080f, 'h103bc, 'h1073f, 'h10794, 'h10747, 'h1074f, 'h10795, 'h10757, 'h106df, 'h10796, 'h10817, 'h106e7, 'h106ef, 'h10797, 'h106f7, 'h106ff, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10799, 'h103bc, 'h10717, 'h1071f, 'h1079a, 'h10727, 'h1072f, 'h1079b, 'h10737, 'h10817, 'h1073f, 'h1079c, 'h10747, 'h1074f, 'h1079d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1079e, 'h1081f, 'h103bc, 'h106e7, 'h106ef, 'h1079f, 'h106f7, 'h106ff, 'h107a0, 'h10707, 'h1070f, 'h107a1, 'h10717, 'h1071f, 'h107a2, 'h10727, 'h1072f, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1081f, 'h103bc, 'h1073f, 'h107a4, 'h10747, 'h1074f, 'h107a5, 'h10757, 'h106df, 'h107a6, 'h10827, 'h106e7, 'h106ef, 'h107a7, 'h106f7, 'h106ff, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107a9, 'h103bc, 'h10717, 'h1071f, 'h107aa, 'h10727, 'h1072f, 'h107ab, 'h10737, 'h10827, 'h1073f, 'h107ac, 'h10747, 'h1074f, 'h107ad, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h107ae, 'h1082f, 'h103bc, 'h106e7, 'h106ef, 'h107af, 'h106f7, 'h106ff, 'h107b0, 'h10707, 'h1070f, 'h107b1, 'h10717, 'h1071f, 'h107b2, 'h10727, 'h1072f, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1082f, 'h103bc, 'h1073f, 'h107b4, 'h10747, 'h1074f, 'h107b5, 'h10757, 'h106df, 'h107b6, 'h10837, 'h106e7, 'h106ef, 'h107b7, 'h106f7, 'h106ff, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107b9, 'h103bc, 'h10717, 'h1071f, 'h107ba, 'h10727, 'h1072f, 'h107bb, 'h10737, 'h10837, 'h1073f, 'h107bc, 'h10747, 'h1074f, 'h107bd, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h107be, 'h1083f, 'h103bc, 'h106e7, 'h106ef, 'h107bf, 'h106f7, 'h106ff, 'h107c0, 'h10707, 'h1070f, 'h107c1, 'h10717, 'h1071f, 'h107c2, 'h10727, 'h1072f, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1083f, 'h103bc, 'h1073f, 'h107c4, 'h10747, 'h1074f, 'h107c5, 'h10757, 'h106df, 'h107c6, 'h10847, 'h106e7, 'h106ef, 'h107c7, 'h106f7, 'h106ff, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107c9, 'h103bc, 'h10717, 'h1071f, 'h107ca, 'h10727, 'h1072f, 'h107cb, 'h10737, 'h10847, 'h1073f, 'h107cc, 'h10747, 'h1074f, 'h107cd, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h107ce, 'h1084f, 'h103bc, 'h106e7, 'h106ef, 'h107cf, 'h106f7, 'h106ff, 'h107d0, 'h10707, 'h1070f, 'h107d1, 'h10717, 'h1071f, 'h107d2, 'h10727, 'h1072f, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1084f, 'h103bc, 'h1073f, 'h107d4, 'h10747, 'h1074f, 'h107d5, 'h10757, 'h106df, 'h107d6, 'h10857, 'h106e7, 'h106ef, 'h107d7, 'h106f7, 'h106ff, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107d9, 'h103bc, 'h10717, 'h1071f, 'h107da, 'h10727, 'h1072f, 'h107db, 'h10737, 'h10857, 'h1073f, 'h107dc, 'h10747, 'h1074f, 'h107dd, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1075e, 'h107df, 'h103bc, 'h106e7, 'h106ef, 'h1075f, 'h106f7, 'h106ff, 'h10760, 'h10707, 'h1070f, 'h10761, 'h10717, 'h1071f, 'h10762, 'h10727, 'h1072f, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h107df, 'h103bc, 'h1073f, 'h10764, 'h10747, 'h1074f, 'h10765, 'h10757, 'h106df, 'h10766, 'h107e7, 'h106e7, 'h106ef, 'h10767, 'h106f7, 'h106ff, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10769, 'h103bc, 'h10717, 'h1071f, 'h1076a, 'h10727, 'h1072f, 'h1076b, 'h10737, 'h107e7, 'h1073f, 'h1076c, 'h10747, 'h1074f, 'h1076d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1076e, 'h107ef, 'h103bc, 'h106e7, 'h106ef, 'h1076f, 'h106f7, 'h106ff, 'h10770, 'h10707, 'h1070f, 'h10771, 'h10717, 'h1071f, 'h10772, 'h10727, 'h1072f, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h107ef, 'h103bc, 'h1073f, 'h10774, 'h10747, 'h1074f, 'h10775, 'h10757, 'h106df, 'h10776, 'h107f7, 'h106e7, 'h106ef, 'h10777, 'h106f7, 'h106ff, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10779, 'h103bc, 'h10717, 'h1071f, 'h1077a, 'h10727, 'h1072f, 'h1077b, 'h10737, 'h107f7, 'h1073f, 'h1077c, 'h10747, 'h1074f, 'h1077d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1077e, 'h107ff, 'h103bc, 'h106e7, 'h106ef, 'h1077f, 'h106f7, 'h106ff, 'h10780, 'h10707, 'h1070f, 'h10781, 'h10717, 'h1071f, 'h10782, 'h10727, 'h1072f, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h107ff, 'h103bc, 'h1073f, 'h10784, 'h10747, 'h1074f, 'h10785, 'h10757, 'h106df, 'h10786, 'h10807, 'h106e7, 'h106ef, 'h10787, 'h106f7, 'h106ff, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10789, 'h103bc, 'h10717, 'h1071f, 'h1078a, 'h10727, 'h1072f, 'h1078b, 'h10737, 'h10807, 'h1073f, 'h1078c, 'h10747, 'h1074f, 'h1078d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1078e, 'h1080f, 'h103bc, 'h106e7, 'h106ef, 'h1078f, 'h106f7, 'h106ff, 'h10790, 'h10707, 'h1070f, 'h10791, 'h10717, 'h1071f, 'h10792, 'h10727, 'h1072f, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1080f, 'h103bc, 'h1073f, 'h10794, 'h10747, 'h1074f, 'h10795, 'h10757, 'h106df, 'h10796, 'h10817, 'h106e7, 'h106ef, 'h10797, 'h106f7, 'h106ff, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h10799, 'h103bc, 'h10717, 'h1071f, 'h1079a, 'h10727, 'h1072f, 'h1079b, 'h10737, 'h10817, 'h1073f, 'h1079c, 'h10747, 'h1074f, 'h1079d, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h1079e, 'h1081f, 'h103bc, 'h106e7, 'h106ef, 'h1079f, 'h106f7, 'h106ff, 'h107a0, 'h10707, 'h1070f, 'h107a1, 'h10717, 'h1071f, 'h107a2, 'h10727, 'h1072f, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1081f, 'h103bc, 'h1073f, 'h107a4, 'h10747, 'h1074f, 'h107a5, 'h10757, 'h106df, 'h107a6, 'h10827, 'h106e7, 'h106ef, 'h107a7, 'h106f7, 'h106ff, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107a9, 'h103bc, 'h10717, 'h1071f, 'h107aa, 'h10727, 'h1072f, 'h107ab, 'h10737, 'h10827, 'h1073f, 'h107ac, 'h10747, 'h1074f, 'h107ad, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h107ae, 'h1082f, 'h103bc, 'h106e7, 'h106ef, 'h107af, 'h106f7, 'h106ff, 'h107b0, 'h10707, 'h1070f, 'h107b1, 'h10717, 'h1071f, 'h107b2, 'h10727, 'h1072f, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1082f, 'h103bc, 'h1073f, 'h107b4, 'h10747, 'h1074f, 'h107b5, 'h10757, 'h106df, 'h107b6, 'h10837, 'h106e7, 'h106ef, 'h107b7, 'h106f7, 'h106ff, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107b9, 'h103bc, 'h10717, 'h1071f, 'h107ba, 'h10727, 'h1072f, 'h107bb, 'h10737, 'h10837, 'h1073f, 'h107bc, 'h10747, 'h1074f, 'h107bd, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h107be, 'h1083f, 'h103bc, 'h106e7, 'h106ef, 'h107bf, 'h106f7, 'h106ff, 'h107c0, 'h10707, 'h1070f, 'h107c1, 'h10717, 'h1071f, 'h107c2, 'h10727, 'h1072f, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1083f, 'h103bc, 'h1073f, 'h107c4, 'h10747, 'h1074f, 'h107c5, 'h10757, 'h106df, 'h107c6, 'h10847, 'h106e7, 'h106ef, 'h107c7, 'h106f7, 'h106ff, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107c9, 'h103bc, 'h10717, 'h1071f, 'h107ca, 'h10727, 'h1072f, 'h107cb, 'h10737, 'h10847, 'h1073f, 'h107cc, 'h10747, 'h1074f, 'h107cd, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106df, 'h107ce, 'h1084f, 'h103bc, 'h106e7, 'h106ef, 'h107cf, 'h106f7, 'h106ff, 'h107d0, 'h10707, 'h1070f, 'h107d1, 'h10717, 'h1071f, 'h107d2, 'h10727, 'h1072f, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h1084f, 'h103bc, 'h1073f, 'h107d4, 'h10747, 'h1074f, 'h107d5, 'h10757, 'h106df, 'h107d6, 'h10857, 'h106e7, 'h106ef, 'h107d7, 'h106f7, 'h106ff, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1070f, 'h107d9, 'h103bc, 'h10717, 'h1071f, 'h107da, 'h10727, 'h1072f, 'h107db, 'h10737, 'h10857, 'h1073f, 'h107dc, 'h10747, 'h1074f, 'h107dd, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1075e, 'h107e0, 'h103bc, 'h106e8, 'h106f0, 'h1075f, 'h106f8, 'h10700, 'h10760, 'h10708, 'h10710, 'h10761, 'h10718, 'h10720, 'h10762, 'h10728, 'h10730, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h107e0, 'h103bc, 'h10740, 'h10764, 'h10748, 'h10750, 'h10765, 'h10758, 'h106e0, 'h10766, 'h107e8, 'h106e8, 'h106f0, 'h10767, 'h106f8, 'h10700, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10769, 'h103bc, 'h10718, 'h10720, 'h1076a, 'h10728, 'h10730, 'h1076b, 'h10738, 'h107e8, 'h10740, 'h1076c, 'h10748, 'h10750, 'h1076d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1076e, 'h107f0, 'h103bc, 'h106e8, 'h106f0, 'h1076f, 'h106f8, 'h10700, 'h10770, 'h10708, 'h10710, 'h10771, 'h10718, 'h10720, 'h10772, 'h10728, 'h10730, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h107f0, 'h103bc, 'h10740, 'h10774, 'h10748, 'h10750, 'h10775, 'h10758, 'h106e0, 'h10776, 'h107f8, 'h106e8, 'h106f0, 'h10777, 'h106f8, 'h10700, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10779, 'h103bc, 'h10718, 'h10720, 'h1077a, 'h10728, 'h10730, 'h1077b, 'h10738, 'h107f8, 'h10740, 'h1077c, 'h10748, 'h10750, 'h1077d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1077e, 'h10800, 'h103bc, 'h106e8, 'h106f0, 'h1077f, 'h106f8, 'h10700, 'h10780, 'h10708, 'h10710, 'h10781, 'h10718, 'h10720, 'h10782, 'h10728, 'h10730, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10800, 'h103bc, 'h10740, 'h10784, 'h10748, 'h10750, 'h10785, 'h10758, 'h106e0, 'h10786, 'h10808, 'h106e8, 'h106f0, 'h10787, 'h106f8, 'h10700, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10789, 'h103bc, 'h10718, 'h10720, 'h1078a, 'h10728, 'h10730, 'h1078b, 'h10738, 'h10808, 'h10740, 'h1078c, 'h10748, 'h10750, 'h1078d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1078e, 'h10810, 'h103bc, 'h106e8, 'h106f0, 'h1078f, 'h106f8, 'h10700, 'h10790, 'h10708, 'h10710, 'h10791, 'h10718, 'h10720, 'h10792, 'h10728, 'h10730, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10810, 'h103bc, 'h10740, 'h10794, 'h10748, 'h10750, 'h10795, 'h10758, 'h106e0, 'h10796, 'h10818, 'h106e8, 'h106f0, 'h10797, 'h106f8, 'h10700, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10799, 'h103bc, 'h10718, 'h10720, 'h1079a, 'h10728, 'h10730, 'h1079b, 'h10738, 'h10818, 'h10740, 'h1079c, 'h10748, 'h10750, 'h1079d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1079e, 'h10820, 'h103bc, 'h106e8, 'h106f0, 'h1079f, 'h106f8, 'h10700, 'h107a0, 'h10708, 'h10710, 'h107a1, 'h10718, 'h10720, 'h107a2, 'h10728, 'h10730, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10820, 'h103bc, 'h10740, 'h107a4, 'h10748, 'h10750, 'h107a5, 'h10758, 'h106e0, 'h107a6, 'h10828, 'h106e8, 'h106f0, 'h107a7, 'h106f8, 'h10700, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107a9, 'h103bc, 'h10718, 'h10720, 'h107aa, 'h10728, 'h10730, 'h107ab, 'h10738, 'h10828, 'h10740, 'h107ac, 'h10748, 'h10750, 'h107ad, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h107ae, 'h10830, 'h103bc, 'h106e8, 'h106f0, 'h107af, 'h106f8, 'h10700, 'h107b0, 'h10708, 'h10710, 'h107b1, 'h10718, 'h10720, 'h107b2, 'h10728, 'h10730, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10830, 'h103bc, 'h10740, 'h107b4, 'h10748, 'h10750, 'h107b5, 'h10758, 'h106e0, 'h107b6, 'h10838, 'h106e8, 'h106f0, 'h107b7, 'h106f8, 'h10700, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107b9, 'h103bc, 'h10718, 'h10720, 'h107ba, 'h10728, 'h10730, 'h107bb, 'h10738, 'h10838, 'h10740, 'h107bc, 'h10748, 'h10750, 'h107bd, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h107be, 'h10840, 'h103bc, 'h106e8, 'h106f0, 'h107bf, 'h106f8, 'h10700, 'h107c0, 'h10708, 'h10710, 'h107c1, 'h10718, 'h10720, 'h107c2, 'h10728, 'h10730, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10840, 'h103bc, 'h10740, 'h107c4, 'h10748, 'h10750, 'h107c5, 'h10758, 'h106e0, 'h107c6, 'h10848, 'h106e8, 'h106f0, 'h107c7, 'h106f8, 'h10700, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107c9, 'h103bc, 'h10718, 'h10720, 'h107ca, 'h10728, 'h10730, 'h107cb, 'h10738, 'h10848, 'h10740, 'h107cc, 'h10748, 'h10750, 'h107cd, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h107ce, 'h10850, 'h103bc, 'h106e8, 'h106f0, 'h107cf, 'h106f8, 'h10700, 'h107d0, 'h10708, 'h10710, 'h107d1, 'h10718, 'h10720, 'h107d2, 'h10728, 'h10730, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10850, 'h103bc, 'h10740, 'h107d4, 'h10748, 'h10750, 'h107d5, 'h10758, 'h106e0, 'h107d6, 'h10858, 'h106e8, 'h106f0, 'h107d7, 'h106f8, 'h10700, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107d9, 'h103bc, 'h10718, 'h10720, 'h107da, 'h10728, 'h10730, 'h107db, 'h10738, 'h10858, 'h10740, 'h107dc, 'h10748, 'h10750, 'h107dd, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1075e, 'h107e0, 'h103bc, 'h106e8, 'h106f0, 'h1075f, 'h106f8, 'h10700, 'h10760, 'h10708, 'h10710, 'h10761, 'h10718, 'h10720, 'h10762, 'h10728, 'h10730, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h107e0, 'h103bc, 'h10740, 'h10764, 'h10748, 'h10750, 'h10765, 'h10758, 'h106e0, 'h10766, 'h107e8, 'h106e8, 'h106f0, 'h10767, 'h106f8, 'h10700, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10769, 'h103bc, 'h10718, 'h10720, 'h1076a, 'h10728, 'h10730, 'h1076b, 'h10738, 'h107e8, 'h10740, 'h1076c, 'h10748, 'h10750, 'h1076d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1076e, 'h107f0, 'h103bc, 'h106e8, 'h106f0, 'h1076f, 'h106f8, 'h10700, 'h10770, 'h10708, 'h10710, 'h10771, 'h10718, 'h10720, 'h10772, 'h10728, 'h10730, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h107f0, 'h103bc, 'h10740, 'h10774, 'h10748, 'h10750, 'h10775, 'h10758, 'h106e0, 'h10776, 'h107f8, 'h106e8, 'h106f0, 'h10777, 'h106f8, 'h10700, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10779, 'h103bc, 'h10718, 'h10720, 'h1077a, 'h10728, 'h10730, 'h1077b, 'h10738, 'h107f8, 'h10740, 'h1077c, 'h10748, 'h10750, 'h1077d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1077e, 'h10800, 'h103bc, 'h106e8, 'h106f0, 'h1077f, 'h106f8, 'h10700, 'h10780, 'h10708, 'h10710, 'h10781, 'h10718, 'h10720, 'h10782, 'h10728, 'h10730, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10800, 'h103bc, 'h10740, 'h10784, 'h10748, 'h10750, 'h10785, 'h10758, 'h106e0, 'h10786, 'h10808, 'h106e8, 'h106f0, 'h10787, 'h106f8, 'h10700, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10789, 'h103bc, 'h10718, 'h10720, 'h1078a, 'h10728, 'h10730, 'h1078b, 'h10738, 'h10808, 'h10740, 'h1078c, 'h10748, 'h10750, 'h1078d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1078e, 'h10810, 'h103bc, 'h106e8, 'h106f0, 'h1078f, 'h106f8, 'h10700, 'h10790, 'h10708, 'h10710, 'h10791, 'h10718, 'h10720, 'h10792, 'h10728, 'h10730, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10810, 'h103bc, 'h10740, 'h10794, 'h10748, 'h10750, 'h10795, 'h10758, 'h106e0, 'h10796, 'h10818, 'h106e8, 'h106f0, 'h10797, 'h106f8, 'h10700, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h10799, 'h103bc, 'h10718, 'h10720, 'h1079a, 'h10728, 'h10730, 'h1079b, 'h10738, 'h10818, 'h10740, 'h1079c, 'h10748, 'h10750, 'h1079d, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h1079e, 'h10820, 'h103bc, 'h106e8, 'h106f0, 'h1079f, 'h106f8, 'h10700, 'h107a0, 'h10708, 'h10710, 'h107a1, 'h10718, 'h10720, 'h107a2, 'h10728, 'h10730, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10820, 'h103bc, 'h10740, 'h107a4, 'h10748, 'h10750, 'h107a5, 'h10758, 'h106e0, 'h107a6, 'h10828, 'h106e8, 'h106f0, 'h107a7, 'h106f8, 'h10700, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107a9, 'h103bc, 'h10718, 'h10720, 'h107aa, 'h10728, 'h10730, 'h107ab, 'h10738, 'h10828, 'h10740, 'h107ac, 'h10748, 'h10750, 'h107ad, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h107ae, 'h10830, 'h103bc, 'h106e8, 'h106f0, 'h107af, 'h106f8, 'h10700, 'h107b0, 'h10708, 'h10710, 'h107b1, 'h10718, 'h10720, 'h107b2, 'h10728, 'h10730, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10830, 'h103bc, 'h10740, 'h107b4, 'h10748, 'h10750, 'h107b5, 'h10758, 'h106e0, 'h107b6, 'h10838, 'h106e8, 'h106f0, 'h107b7, 'h106f8, 'h10700, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107b9, 'h103bc, 'h10718, 'h10720, 'h107ba, 'h10728, 'h10730, 'h107bb, 'h10738, 'h10838, 'h10740, 'h107bc, 'h10748, 'h10750, 'h107bd, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h107be, 'h10840, 'h103bc, 'h106e8, 'h106f0, 'h107bf, 'h106f8, 'h10700, 'h107c0, 'h10708, 'h10710, 'h107c1, 'h10718, 'h10720, 'h107c2, 'h10728, 'h10730, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10840, 'h103bc, 'h10740, 'h107c4, 'h10748, 'h10750, 'h107c5, 'h10758, 'h106e0, 'h107c6, 'h10848, 'h106e8, 'h106f0, 'h107c7, 'h106f8, 'h10700, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107c9, 'h103bc, 'h10718, 'h10720, 'h107ca, 'h10728, 'h10730, 'h107cb, 'h10738, 'h10848, 'h10740, 'h107cc, 'h10748, 'h10750, 'h107cd, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e0, 'h107ce, 'h10850, 'h103bc, 'h106e8, 'h106f0, 'h107cf, 'h106f8, 'h10700, 'h107d0, 'h10708, 'h10710, 'h107d1, 'h10718, 'h10720, 'h107d2, 'h10728, 'h10730, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10738, 'h10850, 'h103bc, 'h10740, 'h107d4, 'h10748, 'h10750, 'h107d5, 'h10758, 'h106e0, 'h107d6, 'h10858, 'h106e8, 'h106f0, 'h107d7, 'h106f8, 'h10700, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10708, 'h10710, 'h107d9, 'h103bc, 'h10718, 'h10720, 'h107da, 'h10728, 'h10730, 'h107db, 'h10738, 'h10858, 'h10740, 'h107dc, 'h10748, 'h10750, 'h107dd, 'h10758, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1075e, 'h107e1, 'h103bc, 'h106e9, 'h106f1, 'h1075f, 'h106f9, 'h10701, 'h10760, 'h10709, 'h10711, 'h10761, 'h10719, 'h10721, 'h10762, 'h10729, 'h10731, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h107e1, 'h103bc, 'h10741, 'h10764, 'h10749, 'h10751, 'h10765, 'h10759, 'h106e1, 'h10766, 'h107e9, 'h106e9, 'h106f1, 'h10767, 'h106f9, 'h10701, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10769, 'h103bc, 'h10719, 'h10721, 'h1076a, 'h10729, 'h10731, 'h1076b, 'h10739, 'h107e9, 'h10741, 'h1076c, 'h10749, 'h10751, 'h1076d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1076e, 'h107f1, 'h103bc, 'h106e9, 'h106f1, 'h1076f, 'h106f9, 'h10701, 'h10770, 'h10709, 'h10711, 'h10771, 'h10719, 'h10721, 'h10772, 'h10729, 'h10731, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h107f1, 'h103bc, 'h10741, 'h10774, 'h10749, 'h10751, 'h10775, 'h10759, 'h106e1, 'h10776, 'h107f9, 'h106e9, 'h106f1, 'h10777, 'h106f9, 'h10701, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10779, 'h103bc, 'h10719, 'h10721, 'h1077a, 'h10729, 'h10731, 'h1077b, 'h10739, 'h107f9, 'h10741, 'h1077c, 'h10749, 'h10751, 'h1077d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1077e, 'h10801, 'h103bc, 'h106e9, 'h106f1, 'h1077f, 'h106f9, 'h10701, 'h10780, 'h10709, 'h10711, 'h10781, 'h10719, 'h10721, 'h10782, 'h10729, 'h10731, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10801, 'h103bc, 'h10741, 'h10784, 'h10749, 'h10751, 'h10785, 'h10759, 'h106e1, 'h10786, 'h10809, 'h106e9, 'h106f1, 'h10787, 'h106f9, 'h10701, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10789, 'h103bc, 'h10719, 'h10721, 'h1078a, 'h10729, 'h10731, 'h1078b, 'h10739, 'h10809, 'h10741, 'h1078c, 'h10749, 'h10751, 'h1078d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1078e, 'h10811, 'h103bc, 'h106e9, 'h106f1, 'h1078f, 'h106f9, 'h10701, 'h10790, 'h10709, 'h10711, 'h10791, 'h10719, 'h10721, 'h10792, 'h10729, 'h10731, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10811, 'h103bc, 'h10741, 'h10794, 'h10749, 'h10751, 'h10795, 'h10759, 'h106e1, 'h10796, 'h10819, 'h106e9, 'h106f1, 'h10797, 'h106f9, 'h10701, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10799, 'h103bc, 'h10719, 'h10721, 'h1079a, 'h10729, 'h10731, 'h1079b, 'h10739, 'h10819, 'h10741, 'h1079c, 'h10749, 'h10751, 'h1079d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1079e, 'h10821, 'h103bc, 'h106e9, 'h106f1, 'h1079f, 'h106f9, 'h10701, 'h107a0, 'h10709, 'h10711, 'h107a1, 'h10719, 'h10721, 'h107a2, 'h10729, 'h10731, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10821, 'h103bc, 'h10741, 'h107a4, 'h10749, 'h10751, 'h107a5, 'h10759, 'h106e1, 'h107a6, 'h10829, 'h106e9, 'h106f1, 'h107a7, 'h106f9, 'h10701, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107a9, 'h103bc, 'h10719, 'h10721, 'h107aa, 'h10729, 'h10731, 'h107ab, 'h10739, 'h10829, 'h10741, 'h107ac, 'h10749, 'h10751, 'h107ad, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h107ae, 'h10831, 'h103bc, 'h106e9, 'h106f1, 'h107af, 'h106f9, 'h10701, 'h107b0, 'h10709, 'h10711, 'h107b1, 'h10719, 'h10721, 'h107b2, 'h10729, 'h10731, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10831, 'h103bc, 'h10741, 'h107b4, 'h10749, 'h10751, 'h107b5, 'h10759, 'h106e1, 'h107b6, 'h10839, 'h106e9, 'h106f1, 'h107b7, 'h106f9, 'h10701, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107b9, 'h103bc, 'h10719, 'h10721, 'h107ba, 'h10729, 'h10731, 'h107bb, 'h10739, 'h10839, 'h10741, 'h107bc, 'h10749, 'h10751, 'h107bd, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h107be, 'h10841, 'h103bc, 'h106e9, 'h106f1, 'h107bf, 'h106f9, 'h10701, 'h107c0, 'h10709, 'h10711, 'h107c1, 'h10719, 'h10721, 'h107c2, 'h10729, 'h10731, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10841, 'h103bc, 'h10741, 'h107c4, 'h10749, 'h10751, 'h107c5, 'h10759, 'h106e1, 'h107c6, 'h10849, 'h106e9, 'h106f1, 'h107c7, 'h106f9, 'h10701, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107c9, 'h103bc, 'h10719, 'h10721, 'h107ca, 'h10729, 'h10731, 'h107cb, 'h10739, 'h10849, 'h10741, 'h107cc, 'h10749, 'h10751, 'h107cd, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h107ce, 'h10851, 'h103bc, 'h106e9, 'h106f1, 'h107cf, 'h106f9, 'h10701, 'h107d0, 'h10709, 'h10711, 'h107d1, 'h10719, 'h10721, 'h107d2, 'h10729, 'h10731, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10851, 'h103bc, 'h10741, 'h107d4, 'h10749, 'h10751, 'h107d5, 'h10759, 'h106e1, 'h107d6, 'h10859, 'h106e9, 'h106f1, 'h107d7, 'h106f9, 'h10701, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107d9, 'h103bc, 'h10719, 'h10721, 'h107da, 'h10729, 'h10731, 'h107db, 'h10739, 'h10859, 'h10741, 'h107dc, 'h10749, 'h10751, 'h107dd, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1075e, 'h107e1, 'h103bc, 'h106e9, 'h106f1, 'h1075f, 'h106f9, 'h10701, 'h10760, 'h10709, 'h10711, 'h10761, 'h10719, 'h10721, 'h10762, 'h10729, 'h10731, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h107e1, 'h103bc, 'h10741, 'h10764, 'h10749, 'h10751, 'h10765, 'h10759, 'h106e1, 'h10766, 'h107e9, 'h106e9, 'h106f1, 'h10767, 'h106f9, 'h10701, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10769, 'h103bc, 'h10719, 'h10721, 'h1076a, 'h10729, 'h10731, 'h1076b, 'h10739, 'h107e9, 'h10741, 'h1076c, 'h10749, 'h10751, 'h1076d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1076e, 'h107f1, 'h103bc, 'h106e9, 'h106f1, 'h1076f, 'h106f9, 'h10701, 'h10770, 'h10709, 'h10711, 'h10771, 'h10719, 'h10721, 'h10772, 'h10729, 'h10731, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h107f1, 'h103bc, 'h10741, 'h10774, 'h10749, 'h10751, 'h10775, 'h10759, 'h106e1, 'h10776, 'h107f9, 'h106e9, 'h106f1, 'h10777, 'h106f9, 'h10701, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10779, 'h103bc, 'h10719, 'h10721, 'h1077a, 'h10729, 'h10731, 'h1077b, 'h10739, 'h107f9, 'h10741, 'h1077c, 'h10749, 'h10751, 'h1077d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1077e, 'h10801, 'h103bc, 'h106e9, 'h106f1, 'h1077f, 'h106f9, 'h10701, 'h10780, 'h10709, 'h10711, 'h10781, 'h10719, 'h10721, 'h10782, 'h10729, 'h10731, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10801, 'h103bc, 'h10741, 'h10784, 'h10749, 'h10751, 'h10785, 'h10759, 'h106e1, 'h10786, 'h10809, 'h106e9, 'h106f1, 'h10787, 'h106f9, 'h10701, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10789, 'h103bc, 'h10719, 'h10721, 'h1078a, 'h10729, 'h10731, 'h1078b, 'h10739, 'h10809, 'h10741, 'h1078c, 'h10749, 'h10751, 'h1078d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1078e, 'h10811, 'h103bc, 'h106e9, 'h106f1, 'h1078f, 'h106f9, 'h10701, 'h10790, 'h10709, 'h10711, 'h10791, 'h10719, 'h10721, 'h10792, 'h10729, 'h10731, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10811, 'h103bc, 'h10741, 'h10794, 'h10749, 'h10751, 'h10795, 'h10759, 'h106e1, 'h10796, 'h10819, 'h106e9, 'h106f1, 'h10797, 'h106f9, 'h10701, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h10799, 'h103bc, 'h10719, 'h10721, 'h1079a, 'h10729, 'h10731, 'h1079b, 'h10739, 'h10819, 'h10741, 'h1079c, 'h10749, 'h10751, 'h1079d, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h1079e, 'h10821, 'h103bc, 'h106e9, 'h106f1, 'h1079f, 'h106f9, 'h10701, 'h107a0, 'h10709, 'h10711, 'h107a1, 'h10719, 'h10721, 'h107a2, 'h10729, 'h10731, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10821, 'h103bc, 'h10741, 'h107a4, 'h10749, 'h10751, 'h107a5, 'h10759, 'h106e1, 'h107a6, 'h10829, 'h106e9, 'h106f1, 'h107a7, 'h106f9, 'h10701, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107a9, 'h103bc, 'h10719, 'h10721, 'h107aa, 'h10729, 'h10731, 'h107ab, 'h10739, 'h10829, 'h10741, 'h107ac, 'h10749, 'h10751, 'h107ad, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h107ae, 'h10831, 'h103bc, 'h106e9, 'h106f1, 'h107af, 'h106f9, 'h10701, 'h107b0, 'h10709, 'h10711, 'h107b1, 'h10719, 'h10721, 'h107b2, 'h10729, 'h10731, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10831, 'h103bc, 'h10741, 'h107b4, 'h10749, 'h10751, 'h107b5, 'h10759, 'h106e1, 'h107b6, 'h10839, 'h106e9, 'h106f1, 'h107b7, 'h106f9, 'h10701, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107b9, 'h103bc, 'h10719, 'h10721, 'h107ba, 'h10729, 'h10731, 'h107bb, 'h10739, 'h10839, 'h10741, 'h107bc, 'h10749, 'h10751, 'h107bd, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h107be, 'h10841, 'h103bc, 'h106e9, 'h106f1, 'h107bf, 'h106f9, 'h10701, 'h107c0, 'h10709, 'h10711, 'h107c1, 'h10719, 'h10721, 'h107c2, 'h10729, 'h10731, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10841, 'h103bc, 'h10741, 'h107c4, 'h10749, 'h10751, 'h107c5, 'h10759, 'h106e1, 'h107c6, 'h10849, 'h106e9, 'h106f1, 'h107c7, 'h106f9, 'h10701, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107c9, 'h103bc, 'h10719, 'h10721, 'h107ca, 'h10729, 'h10731, 'h107cb, 'h10739, 'h10849, 'h10741, 'h107cc, 'h10749, 'h10751, 'h107cd, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e1, 'h107ce, 'h10851, 'h103bc, 'h106e9, 'h106f1, 'h107cf, 'h106f9, 'h10701, 'h107d0, 'h10709, 'h10711, 'h107d1, 'h10719, 'h10721, 'h107d2, 'h10729, 'h10731, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10739, 'h10851, 'h103bc, 'h10741, 'h107d4, 'h10749, 'h10751, 'h107d5, 'h10759, 'h106e1, 'h107d6, 'h10859, 'h106e9, 'h106f1, 'h107d7, 'h106f9, 'h10701, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10709, 'h10711, 'h107d9, 'h103bc, 'h10719, 'h10721, 'h107da, 'h10729, 'h10731, 'h107db, 'h10739, 'h10859, 'h10741, 'h107dc, 'h10749, 'h10751, 'h107dd, 'h10759, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1075e, 'h107e2, 'h103bc, 'h106ea, 'h106f2, 'h1075f, 'h106fa, 'h10702, 'h10760, 'h1070a, 'h10712, 'h10761, 'h1071a, 'h10722, 'h10762, 'h1072a, 'h10732, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h107e2, 'h103bc, 'h10742, 'h10764, 'h1074a, 'h10752, 'h10765, 'h1075a, 'h106e2, 'h10766, 'h107ea, 'h106ea, 'h106f2, 'h10767, 'h106fa, 'h10702, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10769, 'h103bc, 'h1071a, 'h10722, 'h1076a, 'h1072a, 'h10732, 'h1076b, 'h1073a, 'h107ea, 'h10742, 'h1076c, 'h1074a, 'h10752, 'h1076d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1076e, 'h107f2, 'h103bc, 'h106ea, 'h106f2, 'h1076f, 'h106fa, 'h10702, 'h10770, 'h1070a, 'h10712, 'h10771, 'h1071a, 'h10722, 'h10772, 'h1072a, 'h10732, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h107f2, 'h103bc, 'h10742, 'h10774, 'h1074a, 'h10752, 'h10775, 'h1075a, 'h106e2, 'h10776, 'h107fa, 'h106ea, 'h106f2, 'h10777, 'h106fa, 'h10702, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10779, 'h103bc, 'h1071a, 'h10722, 'h1077a, 'h1072a, 'h10732, 'h1077b, 'h1073a, 'h107fa, 'h10742, 'h1077c, 'h1074a, 'h10752, 'h1077d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1077e, 'h10802, 'h103bc, 'h106ea, 'h106f2, 'h1077f, 'h106fa, 'h10702, 'h10780, 'h1070a, 'h10712, 'h10781, 'h1071a, 'h10722, 'h10782, 'h1072a, 'h10732, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10802, 'h103bc, 'h10742, 'h10784, 'h1074a, 'h10752, 'h10785, 'h1075a, 'h106e2, 'h10786, 'h1080a, 'h106ea, 'h106f2, 'h10787, 'h106fa, 'h10702, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10789, 'h103bc, 'h1071a, 'h10722, 'h1078a, 'h1072a, 'h10732, 'h1078b, 'h1073a, 'h1080a, 'h10742, 'h1078c, 'h1074a, 'h10752, 'h1078d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1078e, 'h10812, 'h103bc, 'h106ea, 'h106f2, 'h1078f, 'h106fa, 'h10702, 'h10790, 'h1070a, 'h10712, 'h10791, 'h1071a, 'h10722, 'h10792, 'h1072a, 'h10732, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10812, 'h103bc, 'h10742, 'h10794, 'h1074a, 'h10752, 'h10795, 'h1075a, 'h106e2, 'h10796, 'h1081a, 'h106ea, 'h106f2, 'h10797, 'h106fa, 'h10702, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10799, 'h103bc, 'h1071a, 'h10722, 'h1079a, 'h1072a, 'h10732, 'h1079b, 'h1073a, 'h1081a, 'h10742, 'h1079c, 'h1074a, 'h10752, 'h1079d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1079e, 'h10822, 'h103bc, 'h106ea, 'h106f2, 'h1079f, 'h106fa, 'h10702, 'h107a0, 'h1070a, 'h10712, 'h107a1, 'h1071a, 'h10722, 'h107a2, 'h1072a, 'h10732, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10822, 'h103bc, 'h10742, 'h107a4, 'h1074a, 'h10752, 'h107a5, 'h1075a, 'h106e2, 'h107a6, 'h1082a, 'h106ea, 'h106f2, 'h107a7, 'h106fa, 'h10702, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107a9, 'h103bc, 'h1071a, 'h10722, 'h107aa, 'h1072a, 'h10732, 'h107ab, 'h1073a, 'h1082a, 'h10742, 'h107ac, 'h1074a, 'h10752, 'h107ad, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h107ae, 'h10832, 'h103bc, 'h106ea, 'h106f2, 'h107af, 'h106fa, 'h10702, 'h107b0, 'h1070a, 'h10712, 'h107b1, 'h1071a, 'h10722, 'h107b2, 'h1072a, 'h10732, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10832, 'h103bc, 'h10742, 'h107b4, 'h1074a, 'h10752, 'h107b5, 'h1075a, 'h106e2, 'h107b6, 'h1083a, 'h106ea, 'h106f2, 'h107b7, 'h106fa, 'h10702, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107b9, 'h103bc, 'h1071a, 'h10722, 'h107ba, 'h1072a, 'h10732, 'h107bb, 'h1073a, 'h1083a, 'h10742, 'h107bc, 'h1074a, 'h10752, 'h107bd, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h107be, 'h10842, 'h103bc, 'h106ea, 'h106f2, 'h107bf, 'h106fa, 'h10702, 'h107c0, 'h1070a, 'h10712, 'h107c1, 'h1071a, 'h10722, 'h107c2, 'h1072a, 'h10732, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10842, 'h103bc, 'h10742, 'h107c4, 'h1074a, 'h10752, 'h107c5, 'h1075a, 'h106e2, 'h107c6, 'h1084a, 'h106ea, 'h106f2, 'h107c7, 'h106fa, 'h10702, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107c9, 'h103bc, 'h1071a, 'h10722, 'h107ca, 'h1072a, 'h10732, 'h107cb, 'h1073a, 'h1084a, 'h10742, 'h107cc, 'h1074a, 'h10752, 'h107cd, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h107ce, 'h10852, 'h103bc, 'h106ea, 'h106f2, 'h107cf, 'h106fa, 'h10702, 'h107d0, 'h1070a, 'h10712, 'h107d1, 'h1071a, 'h10722, 'h107d2, 'h1072a, 'h10732, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10852, 'h103bc, 'h10742, 'h107d4, 'h1074a, 'h10752, 'h107d5, 'h1075a, 'h106e2, 'h107d6, 'h1085a, 'h106ea, 'h106f2, 'h107d7, 'h106fa, 'h10702, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107d9, 'h103bc, 'h1071a, 'h10722, 'h107da, 'h1072a, 'h10732, 'h107db, 'h1073a, 'h1085a, 'h10742, 'h107dc, 'h1074a, 'h10752, 'h107dd, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1075e, 'h107e2, 'h103bc, 'h106ea, 'h106f2, 'h1075f, 'h106fa, 'h10702, 'h10760, 'h1070a, 'h10712, 'h10761, 'h1071a, 'h10722, 'h10762, 'h1072a, 'h10732, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h107e2, 'h103bc, 'h10742, 'h10764, 'h1074a, 'h10752, 'h10765, 'h1075a, 'h106e2, 'h10766, 'h107ea, 'h106ea, 'h106f2, 'h10767, 'h106fa, 'h10702, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10769, 'h103bc, 'h1071a, 'h10722, 'h1076a, 'h1072a, 'h10732, 'h1076b, 'h1073a, 'h107ea, 'h10742, 'h1076c, 'h1074a, 'h10752, 'h1076d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1076e, 'h107f2, 'h103bc, 'h106ea, 'h106f2, 'h1076f, 'h106fa, 'h10702, 'h10770, 'h1070a, 'h10712, 'h10771, 'h1071a, 'h10722, 'h10772, 'h1072a, 'h10732, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h107f2, 'h103bc, 'h10742, 'h10774, 'h1074a, 'h10752, 'h10775, 'h1075a, 'h106e2, 'h10776, 'h107fa, 'h106ea, 'h106f2, 'h10777, 'h106fa, 'h10702, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10779, 'h103bc, 'h1071a, 'h10722, 'h1077a, 'h1072a, 'h10732, 'h1077b, 'h1073a, 'h107fa, 'h10742, 'h1077c, 'h1074a, 'h10752, 'h1077d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1077e, 'h10802, 'h103bc, 'h106ea, 'h106f2, 'h1077f, 'h106fa, 'h10702, 'h10780, 'h1070a, 'h10712, 'h10781, 'h1071a, 'h10722, 'h10782, 'h1072a, 'h10732, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10802, 'h103bc, 'h10742, 'h10784, 'h1074a, 'h10752, 'h10785, 'h1075a, 'h106e2, 'h10786, 'h1080a, 'h106ea, 'h106f2, 'h10787, 'h106fa, 'h10702, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10789, 'h103bc, 'h1071a, 'h10722, 'h1078a, 'h1072a, 'h10732, 'h1078b, 'h1073a, 'h1080a, 'h10742, 'h1078c, 'h1074a, 'h10752, 'h1078d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1078e, 'h10812, 'h103bc, 'h106ea, 'h106f2, 'h1078f, 'h106fa, 'h10702, 'h10790, 'h1070a, 'h10712, 'h10791, 'h1071a, 'h10722, 'h10792, 'h1072a, 'h10732, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10812, 'h103bc, 'h10742, 'h10794, 'h1074a, 'h10752, 'h10795, 'h1075a, 'h106e2, 'h10796, 'h1081a, 'h106ea, 'h106f2, 'h10797, 'h106fa, 'h10702, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h10799, 'h103bc, 'h1071a, 'h10722, 'h1079a, 'h1072a, 'h10732, 'h1079b, 'h1073a, 'h1081a, 'h10742, 'h1079c, 'h1074a, 'h10752, 'h1079d, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h1079e, 'h10822, 'h103bc, 'h106ea, 'h106f2, 'h1079f, 'h106fa, 'h10702, 'h107a0, 'h1070a, 'h10712, 'h107a1, 'h1071a, 'h10722, 'h107a2, 'h1072a, 'h10732, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10822, 'h103bc, 'h10742, 'h107a4, 'h1074a, 'h10752, 'h107a5, 'h1075a, 'h106e2, 'h107a6, 'h1082a, 'h106ea, 'h106f2, 'h107a7, 'h106fa, 'h10702, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107a9, 'h103bc, 'h1071a, 'h10722, 'h107aa, 'h1072a, 'h10732, 'h107ab, 'h1073a, 'h1082a, 'h10742, 'h107ac, 'h1074a, 'h10752, 'h107ad, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h107ae, 'h10832, 'h103bc, 'h106ea, 'h106f2, 'h107af, 'h106fa, 'h10702, 'h107b0, 'h1070a, 'h10712, 'h107b1, 'h1071a, 'h10722, 'h107b2, 'h1072a, 'h10732, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10832, 'h103bc, 'h10742, 'h107b4, 'h1074a, 'h10752, 'h107b5, 'h1075a, 'h106e2, 'h107b6, 'h1083a, 'h106ea, 'h106f2, 'h107b7, 'h106fa, 'h10702, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107b9, 'h103bc, 'h1071a, 'h10722, 'h107ba, 'h1072a, 'h10732, 'h107bb, 'h1073a, 'h1083a, 'h10742, 'h107bc, 'h1074a, 'h10752, 'h107bd, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h107be, 'h10842, 'h103bc, 'h106ea, 'h106f2, 'h107bf, 'h106fa, 'h10702, 'h107c0, 'h1070a, 'h10712, 'h107c1, 'h1071a, 'h10722, 'h107c2, 'h1072a, 'h10732, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10842, 'h103bc, 'h10742, 'h107c4, 'h1074a, 'h10752, 'h107c5, 'h1075a, 'h106e2, 'h107c6, 'h1084a, 'h106ea, 'h106f2, 'h107c7, 'h106fa, 'h10702, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107c9, 'h103bc, 'h1071a, 'h10722, 'h107ca, 'h1072a, 'h10732, 'h107cb, 'h1073a, 'h1084a, 'h10742, 'h107cc, 'h1074a, 'h10752, 'h107cd, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e2, 'h107ce, 'h10852, 'h103bc, 'h106ea, 'h106f2, 'h107cf, 'h106fa, 'h10702, 'h107d0, 'h1070a, 'h10712, 'h107d1, 'h1071a, 'h10722, 'h107d2, 'h1072a, 'h10732, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073a, 'h10852, 'h103bc, 'h10742, 'h107d4, 'h1074a, 'h10752, 'h107d5, 'h1075a, 'h106e2, 'h107d6, 'h1085a, 'h106ea, 'h106f2, 'h107d7, 'h106fa, 'h10702, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070a, 'h10712, 'h107d9, 'h103bc, 'h1071a, 'h10722, 'h107da, 'h1072a, 'h10732, 'h107db, 'h1073a, 'h1085a, 'h10742, 'h107dc, 'h1074a, 'h10752, 'h107dd, 'h1075a, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1075e, 'h107e3, 'h103bc, 'h106eb, 'h106f3, 'h1075f, 'h106fb, 'h10703, 'h10760, 'h1070b, 'h10713, 'h10761, 'h1071b, 'h10723, 'h10762, 'h1072b, 'h10733, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h107e3, 'h103bc, 'h10743, 'h10764, 'h1074b, 'h10753, 'h10765, 'h1075b, 'h106e3, 'h10766, 'h107eb, 'h106eb, 'h106f3, 'h10767, 'h106fb, 'h10703, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10769, 'h103bc, 'h1071b, 'h10723, 'h1076a, 'h1072b, 'h10733, 'h1076b, 'h1073b, 'h107eb, 'h10743, 'h1076c, 'h1074b, 'h10753, 'h1076d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1076e, 'h107f3, 'h103bc, 'h106eb, 'h106f3, 'h1076f, 'h106fb, 'h10703, 'h10770, 'h1070b, 'h10713, 'h10771, 'h1071b, 'h10723, 'h10772, 'h1072b, 'h10733, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h107f3, 'h103bc, 'h10743, 'h10774, 'h1074b, 'h10753, 'h10775, 'h1075b, 'h106e3, 'h10776, 'h107fb, 'h106eb, 'h106f3, 'h10777, 'h106fb, 'h10703, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10779, 'h103bc, 'h1071b, 'h10723, 'h1077a, 'h1072b, 'h10733, 'h1077b, 'h1073b, 'h107fb, 'h10743, 'h1077c, 'h1074b, 'h10753, 'h1077d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1077e, 'h10803, 'h103bc, 'h106eb, 'h106f3, 'h1077f, 'h106fb, 'h10703, 'h10780, 'h1070b, 'h10713, 'h10781, 'h1071b, 'h10723, 'h10782, 'h1072b, 'h10733, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10803, 'h103bc, 'h10743, 'h10784, 'h1074b, 'h10753, 'h10785, 'h1075b, 'h106e3, 'h10786, 'h1080b, 'h106eb, 'h106f3, 'h10787, 'h106fb, 'h10703, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10789, 'h103bc, 'h1071b, 'h10723, 'h1078a, 'h1072b, 'h10733, 'h1078b, 'h1073b, 'h1080b, 'h10743, 'h1078c, 'h1074b, 'h10753, 'h1078d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1078e, 'h10813, 'h103bc, 'h106eb, 'h106f3, 'h1078f, 'h106fb, 'h10703, 'h10790, 'h1070b, 'h10713, 'h10791, 'h1071b, 'h10723, 'h10792, 'h1072b, 'h10733, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10813, 'h103bc, 'h10743, 'h10794, 'h1074b, 'h10753, 'h10795, 'h1075b, 'h106e3, 'h10796, 'h1081b, 'h106eb, 'h106f3, 'h10797, 'h106fb, 'h10703, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10799, 'h103bc, 'h1071b, 'h10723, 'h1079a, 'h1072b, 'h10733, 'h1079b, 'h1073b, 'h1081b, 'h10743, 'h1079c, 'h1074b, 'h10753, 'h1079d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1079e, 'h10823, 'h103bc, 'h106eb, 'h106f3, 'h1079f, 'h106fb, 'h10703, 'h107a0, 'h1070b, 'h10713, 'h107a1, 'h1071b, 'h10723, 'h107a2, 'h1072b, 'h10733, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10823, 'h103bc, 'h10743, 'h107a4, 'h1074b, 'h10753, 'h107a5, 'h1075b, 'h106e3, 'h107a6, 'h1082b, 'h106eb, 'h106f3, 'h107a7, 'h106fb, 'h10703, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107a9, 'h103bc, 'h1071b, 'h10723, 'h107aa, 'h1072b, 'h10733, 'h107ab, 'h1073b, 'h1082b, 'h10743, 'h107ac, 'h1074b, 'h10753, 'h107ad, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h107ae, 'h10833, 'h103bc, 'h106eb, 'h106f3, 'h107af, 'h106fb, 'h10703, 'h107b0, 'h1070b, 'h10713, 'h107b1, 'h1071b, 'h10723, 'h107b2, 'h1072b, 'h10733, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10833, 'h103bc, 'h10743, 'h107b4, 'h1074b, 'h10753, 'h107b5, 'h1075b, 'h106e3, 'h107b6, 'h1083b, 'h106eb, 'h106f3, 'h107b7, 'h106fb, 'h10703, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107b9, 'h103bc, 'h1071b, 'h10723, 'h107ba, 'h1072b, 'h10733, 'h107bb, 'h1073b, 'h1083b, 'h10743, 'h107bc, 'h1074b, 'h10753, 'h107bd, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h107be, 'h10843, 'h103bc, 'h106eb, 'h106f3, 'h107bf, 'h106fb, 'h10703, 'h107c0, 'h1070b, 'h10713, 'h107c1, 'h1071b, 'h10723, 'h107c2, 'h1072b, 'h10733, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10843, 'h103bc, 'h10743, 'h107c4, 'h1074b, 'h10753, 'h107c5, 'h1075b, 'h106e3, 'h107c6, 'h1084b, 'h106eb, 'h106f3, 'h107c7, 'h106fb, 'h10703, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107c9, 'h103bc, 'h1071b, 'h10723, 'h107ca, 'h1072b, 'h10733, 'h107cb, 'h1073b, 'h1084b, 'h10743, 'h107cc, 'h1074b, 'h10753, 'h107cd, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h107ce, 'h10853, 'h103bc, 'h106eb, 'h106f3, 'h107cf, 'h106fb, 'h10703, 'h107d0, 'h1070b, 'h10713, 'h107d1, 'h1071b, 'h10723, 'h107d2, 'h1072b, 'h10733, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10853, 'h103bc, 'h10743, 'h107d4, 'h1074b, 'h10753, 'h107d5, 'h1075b, 'h106e3, 'h107d6, 'h1085b, 'h106eb, 'h106f3, 'h107d7, 'h106fb, 'h10703, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107d9, 'h103bc, 'h1071b, 'h10723, 'h107da, 'h1072b, 'h10733, 'h107db, 'h1073b, 'h1085b, 'h10743, 'h107dc, 'h1074b, 'h10753, 'h107dd, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1075e, 'h107e3, 'h103bc, 'h106eb, 'h106f3, 'h1075f, 'h106fb, 'h10703, 'h10760, 'h1070b, 'h10713, 'h10761, 'h1071b, 'h10723, 'h10762, 'h1072b, 'h10733, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h107e3, 'h103bc, 'h10743, 'h10764, 'h1074b, 'h10753, 'h10765, 'h1075b, 'h106e3, 'h10766, 'h107eb, 'h106eb, 'h106f3, 'h10767, 'h106fb, 'h10703, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10769, 'h103bc, 'h1071b, 'h10723, 'h1076a, 'h1072b, 'h10733, 'h1076b, 'h1073b, 'h107eb, 'h10743, 'h1076c, 'h1074b, 'h10753, 'h1076d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1076e, 'h107f3, 'h103bc, 'h106eb, 'h106f3, 'h1076f, 'h106fb, 'h10703, 'h10770, 'h1070b, 'h10713, 'h10771, 'h1071b, 'h10723, 'h10772, 'h1072b, 'h10733, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h107f3, 'h103bc, 'h10743, 'h10774, 'h1074b, 'h10753, 'h10775, 'h1075b, 'h106e3, 'h10776, 'h107fb, 'h106eb, 'h106f3, 'h10777, 'h106fb, 'h10703, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10779, 'h103bc, 'h1071b, 'h10723, 'h1077a, 'h1072b, 'h10733, 'h1077b, 'h1073b, 'h107fb, 'h10743, 'h1077c, 'h1074b, 'h10753, 'h1077d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1077e, 'h10803, 'h103bc, 'h106eb, 'h106f3, 'h1077f, 'h106fb, 'h10703, 'h10780, 'h1070b, 'h10713, 'h10781, 'h1071b, 'h10723, 'h10782, 'h1072b, 'h10733, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10803, 'h103bc, 'h10743, 'h10784, 'h1074b, 'h10753, 'h10785, 'h1075b, 'h106e3, 'h10786, 'h1080b, 'h106eb, 'h106f3, 'h10787, 'h106fb, 'h10703, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10789, 'h103bc, 'h1071b, 'h10723, 'h1078a, 'h1072b, 'h10733, 'h1078b, 'h1073b, 'h1080b, 'h10743, 'h1078c, 'h1074b, 'h10753, 'h1078d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1078e, 'h10813, 'h103bc, 'h106eb, 'h106f3, 'h1078f, 'h106fb, 'h10703, 'h10790, 'h1070b, 'h10713, 'h10791, 'h1071b, 'h10723, 'h10792, 'h1072b, 'h10733, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10813, 'h103bc, 'h10743, 'h10794, 'h1074b, 'h10753, 'h10795, 'h1075b, 'h106e3, 'h10796, 'h1081b, 'h106eb, 'h106f3, 'h10797, 'h106fb, 'h10703, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h10799, 'h103bc, 'h1071b, 'h10723, 'h1079a, 'h1072b, 'h10733, 'h1079b, 'h1073b, 'h1081b, 'h10743, 'h1079c, 'h1074b, 'h10753, 'h1079d, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h1079e, 'h10823, 'h103bc, 'h106eb, 'h106f3, 'h1079f, 'h106fb, 'h10703, 'h107a0, 'h1070b, 'h10713, 'h107a1, 'h1071b, 'h10723, 'h107a2, 'h1072b, 'h10733, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10823, 'h103bc, 'h10743, 'h107a4, 'h1074b, 'h10753, 'h107a5, 'h1075b, 'h106e3, 'h107a6, 'h1082b, 'h106eb, 'h106f3, 'h107a7, 'h106fb, 'h10703, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107a9, 'h103bc, 'h1071b, 'h10723, 'h107aa, 'h1072b, 'h10733, 'h107ab, 'h1073b, 'h1082b, 'h10743, 'h107ac, 'h1074b, 'h10753, 'h107ad, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h107ae, 'h10833, 'h103bc, 'h106eb, 'h106f3, 'h107af, 'h106fb, 'h10703, 'h107b0, 'h1070b, 'h10713, 'h107b1, 'h1071b, 'h10723, 'h107b2, 'h1072b, 'h10733, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10833, 'h103bc, 'h10743, 'h107b4, 'h1074b, 'h10753, 'h107b5, 'h1075b, 'h106e3, 'h107b6, 'h1083b, 'h106eb, 'h106f3, 'h107b7, 'h106fb, 'h10703, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107b9, 'h103bc, 'h1071b, 'h10723, 'h107ba, 'h1072b, 'h10733, 'h107bb, 'h1073b, 'h1083b, 'h10743, 'h107bc, 'h1074b, 'h10753, 'h107bd, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h107be, 'h10843, 'h103bc, 'h106eb, 'h106f3, 'h107bf, 'h106fb, 'h10703, 'h107c0, 'h1070b, 'h10713, 'h107c1, 'h1071b, 'h10723, 'h107c2, 'h1072b, 'h10733, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10843, 'h103bc, 'h10743, 'h107c4, 'h1074b, 'h10753, 'h107c5, 'h1075b, 'h106e3, 'h107c6, 'h1084b, 'h106eb, 'h106f3, 'h107c7, 'h106fb, 'h10703, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107c9, 'h103bc, 'h1071b, 'h10723, 'h107ca, 'h1072b, 'h10733, 'h107cb, 'h1073b, 'h1084b, 'h10743, 'h107cc, 'h1074b, 'h10753, 'h107cd, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e3, 'h107ce, 'h10853, 'h103bc, 'h106eb, 'h106f3, 'h107cf, 'h106fb, 'h10703, 'h107d0, 'h1070b, 'h10713, 'h107d1, 'h1071b, 'h10723, 'h107d2, 'h1072b, 'h10733, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073b, 'h10853, 'h103bc, 'h10743, 'h107d4, 'h1074b, 'h10753, 'h107d5, 'h1075b, 'h106e3, 'h107d6, 'h1085b, 'h106eb, 'h106f3, 'h107d7, 'h106fb, 'h10703, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070b, 'h10713, 'h107d9, 'h103bc, 'h1071b, 'h10723, 'h107da, 'h1072b, 'h10733, 'h107db, 'h1073b, 'h1085b, 'h10743, 'h107dc, 'h1074b, 'h10753, 'h107dd, 'h1075b, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1075e, 'h107e4, 'h103bc, 'h106ec, 'h106f4, 'h1075f, 'h106fc, 'h10704, 'h10760, 'h1070c, 'h10714, 'h10761, 'h1071c, 'h10724, 'h10762, 'h1072c, 'h10734, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h107e4, 'h103bc, 'h10744, 'h10764, 'h1074c, 'h10754, 'h10765, 'h1075c, 'h106e4, 'h10766, 'h107ec, 'h106ec, 'h106f4, 'h10767, 'h106fc, 'h10704, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10769, 'h103bc, 'h1071c, 'h10724, 'h1076a, 'h1072c, 'h10734, 'h1076b, 'h1073c, 'h107ec, 'h10744, 'h1076c, 'h1074c, 'h10754, 'h1076d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1076e, 'h107f4, 'h103bc, 'h106ec, 'h106f4, 'h1076f, 'h106fc, 'h10704, 'h10770, 'h1070c, 'h10714, 'h10771, 'h1071c, 'h10724, 'h10772, 'h1072c, 'h10734, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h107f4, 'h103bc, 'h10744, 'h10774, 'h1074c, 'h10754, 'h10775, 'h1075c, 'h106e4, 'h10776, 'h107fc, 'h106ec, 'h106f4, 'h10777, 'h106fc, 'h10704, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10779, 'h103bc, 'h1071c, 'h10724, 'h1077a, 'h1072c, 'h10734, 'h1077b, 'h1073c, 'h107fc, 'h10744, 'h1077c, 'h1074c, 'h10754, 'h1077d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1077e, 'h10804, 'h103bc, 'h106ec, 'h106f4, 'h1077f, 'h106fc, 'h10704, 'h10780, 'h1070c, 'h10714, 'h10781, 'h1071c, 'h10724, 'h10782, 'h1072c, 'h10734, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10804, 'h103bc, 'h10744, 'h10784, 'h1074c, 'h10754, 'h10785, 'h1075c, 'h106e4, 'h10786, 'h1080c, 'h106ec, 'h106f4, 'h10787, 'h106fc, 'h10704, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10789, 'h103bc, 'h1071c, 'h10724, 'h1078a, 'h1072c, 'h10734, 'h1078b, 'h1073c, 'h1080c, 'h10744, 'h1078c, 'h1074c, 'h10754, 'h1078d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1078e, 'h10814, 'h103bc, 'h106ec, 'h106f4, 'h1078f, 'h106fc, 'h10704, 'h10790, 'h1070c, 'h10714, 'h10791, 'h1071c, 'h10724, 'h10792, 'h1072c, 'h10734, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10814, 'h103bc, 'h10744, 'h10794, 'h1074c, 'h10754, 'h10795, 'h1075c, 'h106e4, 'h10796, 'h1081c, 'h106ec, 'h106f4, 'h10797, 'h106fc, 'h10704, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10799, 'h103bc, 'h1071c, 'h10724, 'h1079a, 'h1072c, 'h10734, 'h1079b, 'h1073c, 'h1081c, 'h10744, 'h1079c, 'h1074c, 'h10754, 'h1079d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1079e, 'h10824, 'h103bc, 'h106ec, 'h106f4, 'h1079f, 'h106fc, 'h10704, 'h107a0, 'h1070c, 'h10714, 'h107a1, 'h1071c, 'h10724, 'h107a2, 'h1072c, 'h10734, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10824, 'h103bc, 'h10744, 'h107a4, 'h1074c, 'h10754, 'h107a5, 'h1075c, 'h106e4, 'h107a6, 'h1082c, 'h106ec, 'h106f4, 'h107a7, 'h106fc, 'h10704, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107a9, 'h103bc, 'h1071c, 'h10724, 'h107aa, 'h1072c, 'h10734, 'h107ab, 'h1073c, 'h1082c, 'h10744, 'h107ac, 'h1074c, 'h10754, 'h107ad, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h107ae, 'h10834, 'h103bc, 'h106ec, 'h106f4, 'h107af, 'h106fc, 'h10704, 'h107b0, 'h1070c, 'h10714, 'h107b1, 'h1071c, 'h10724, 'h107b2, 'h1072c, 'h10734, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10834, 'h103bc, 'h10744, 'h107b4, 'h1074c, 'h10754, 'h107b5, 'h1075c, 'h106e4, 'h107b6, 'h1083c, 'h106ec, 'h106f4, 'h107b7, 'h106fc, 'h10704, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107b9, 'h103bc, 'h1071c, 'h10724, 'h107ba, 'h1072c, 'h10734, 'h107bb, 'h1073c, 'h1083c, 'h10744, 'h107bc, 'h1074c, 'h10754, 'h107bd, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h107be, 'h10844, 'h103bc, 'h106ec, 'h106f4, 'h107bf, 'h106fc, 'h10704, 'h107c0, 'h1070c, 'h10714, 'h107c1, 'h1071c, 'h10724, 'h107c2, 'h1072c, 'h10734, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10844, 'h103bc, 'h10744, 'h107c4, 'h1074c, 'h10754, 'h107c5, 'h1075c, 'h106e4, 'h107c6, 'h1084c, 'h106ec, 'h106f4, 'h107c7, 'h106fc, 'h10704, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107c9, 'h103bc, 'h1071c, 'h10724, 'h107ca, 'h1072c, 'h10734, 'h107cb, 'h1073c, 'h1084c, 'h10744, 'h107cc, 'h1074c, 'h10754, 'h107cd, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h107ce, 'h10854, 'h103bc, 'h106ec, 'h106f4, 'h107cf, 'h106fc, 'h10704, 'h107d0, 'h1070c, 'h10714, 'h107d1, 'h1071c, 'h10724, 'h107d2, 'h1072c, 'h10734, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10854, 'h103bc, 'h10744, 'h107d4, 'h1074c, 'h10754, 'h107d5, 'h1075c, 'h106e4, 'h107d6, 'h1085c, 'h106ec, 'h106f4, 'h107d7, 'h106fc, 'h10704, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107d9, 'h103bc, 'h1071c, 'h10724, 'h107da, 'h1072c, 'h10734, 'h107db, 'h1073c, 'h1085c, 'h10744, 'h107dc, 'h1074c, 'h10754, 'h107dd, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1075e, 'h107e4, 'h103bc, 'h106ec, 'h106f4, 'h1075f, 'h106fc, 'h10704, 'h10760, 'h1070c, 'h10714, 'h10761, 'h1071c, 'h10724, 'h10762, 'h1072c, 'h10734, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h107e4, 'h103bc, 'h10744, 'h10764, 'h1074c, 'h10754, 'h10765, 'h1075c, 'h106e4, 'h10766, 'h107ec, 'h106ec, 'h106f4, 'h10767, 'h106fc, 'h10704, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10769, 'h103bc, 'h1071c, 'h10724, 'h1076a, 'h1072c, 'h10734, 'h1076b, 'h1073c, 'h107ec, 'h10744, 'h1076c, 'h1074c, 'h10754, 'h1076d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1076e, 'h107f4, 'h103bc, 'h106ec, 'h106f4, 'h1076f, 'h106fc, 'h10704, 'h10770, 'h1070c, 'h10714, 'h10771, 'h1071c, 'h10724, 'h10772, 'h1072c, 'h10734, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h107f4, 'h103bc, 'h10744, 'h10774, 'h1074c, 'h10754, 'h10775, 'h1075c, 'h106e4, 'h10776, 'h107fc, 'h106ec, 'h106f4, 'h10777, 'h106fc, 'h10704, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10779, 'h103bc, 'h1071c, 'h10724, 'h1077a, 'h1072c, 'h10734, 'h1077b, 'h1073c, 'h107fc, 'h10744, 'h1077c, 'h1074c, 'h10754, 'h1077d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1077e, 'h10804, 'h103bc, 'h106ec, 'h106f4, 'h1077f, 'h106fc, 'h10704, 'h10780, 'h1070c, 'h10714, 'h10781, 'h1071c, 'h10724, 'h10782, 'h1072c, 'h10734, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10804, 'h103bc, 'h10744, 'h10784, 'h1074c, 'h10754, 'h10785, 'h1075c, 'h106e4, 'h10786, 'h1080c, 'h106ec, 'h106f4, 'h10787, 'h106fc, 'h10704, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10789, 'h103bc, 'h1071c, 'h10724, 'h1078a, 'h1072c, 'h10734, 'h1078b, 'h1073c, 'h1080c, 'h10744, 'h1078c, 'h1074c, 'h10754, 'h1078d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1078e, 'h10814, 'h103bc, 'h106ec, 'h106f4, 'h1078f, 'h106fc, 'h10704, 'h10790, 'h1070c, 'h10714, 'h10791, 'h1071c, 'h10724, 'h10792, 'h1072c, 'h10734, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10814, 'h103bc, 'h10744, 'h10794, 'h1074c, 'h10754, 'h10795, 'h1075c, 'h106e4, 'h10796, 'h1081c, 'h106ec, 'h106f4, 'h10797, 'h106fc, 'h10704, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h10799, 'h103bc, 'h1071c, 'h10724, 'h1079a, 'h1072c, 'h10734, 'h1079b, 'h1073c, 'h1081c, 'h10744, 'h1079c, 'h1074c, 'h10754, 'h1079d, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h1079e, 'h10824, 'h103bc, 'h106ec, 'h106f4, 'h1079f, 'h106fc, 'h10704, 'h107a0, 'h1070c, 'h10714, 'h107a1, 'h1071c, 'h10724, 'h107a2, 'h1072c, 'h10734, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10824, 'h103bc, 'h10744, 'h107a4, 'h1074c, 'h10754, 'h107a5, 'h1075c, 'h106e4, 'h107a6, 'h1082c, 'h106ec, 'h106f4, 'h107a7, 'h106fc, 'h10704, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107a9, 'h103bc, 'h1071c, 'h10724, 'h107aa, 'h1072c, 'h10734, 'h107ab, 'h1073c, 'h1082c, 'h10744, 'h107ac, 'h1074c, 'h10754, 'h107ad, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h107ae, 'h10834, 'h103bc, 'h106ec, 'h106f4, 'h107af, 'h106fc, 'h10704, 'h107b0, 'h1070c, 'h10714, 'h107b1, 'h1071c, 'h10724, 'h107b2, 'h1072c, 'h10734, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10834, 'h103bc, 'h10744, 'h107b4, 'h1074c, 'h10754, 'h107b5, 'h1075c, 'h106e4, 'h107b6, 'h1083c, 'h106ec, 'h106f4, 'h107b7, 'h106fc, 'h10704, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107b9, 'h103bc, 'h1071c, 'h10724, 'h107ba, 'h1072c, 'h10734, 'h107bb, 'h1073c, 'h1083c, 'h10744, 'h107bc, 'h1074c, 'h10754, 'h107bd, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h107be, 'h10844, 'h103bc, 'h106ec, 'h106f4, 'h107bf, 'h106fc, 'h10704, 'h107c0, 'h1070c, 'h10714, 'h107c1, 'h1071c, 'h10724, 'h107c2, 'h1072c, 'h10734, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10844, 'h103bc, 'h10744, 'h107c4, 'h1074c, 'h10754, 'h107c5, 'h1075c, 'h106e4, 'h107c6, 'h1084c, 'h106ec, 'h106f4, 'h107c7, 'h106fc, 'h10704, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107c9, 'h103bc, 'h1071c, 'h10724, 'h107ca, 'h1072c, 'h10734, 'h107cb, 'h1073c, 'h1084c, 'h10744, 'h107cc, 'h1074c, 'h10754, 'h107cd, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e4, 'h107ce, 'h10854, 'h103bc, 'h106ec, 'h106f4, 'h107cf, 'h106fc, 'h10704, 'h107d0, 'h1070c, 'h10714, 'h107d1, 'h1071c, 'h10724, 'h107d2, 'h1072c, 'h10734, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073c, 'h10854, 'h103bc, 'h10744, 'h107d4, 'h1074c, 'h10754, 'h107d5, 'h1075c, 'h106e4, 'h107d6, 'h1085c, 'h106ec, 'h106f4, 'h107d7, 'h106fc, 'h10704, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070c, 'h10714, 'h107d9, 'h103bc, 'h1071c, 'h10724, 'h107da, 'h1072c, 'h10734, 'h107db, 'h1073c, 'h1085c, 'h10744, 'h107dc, 'h1074c, 'h10754, 'h107dd, 'h1075c, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1075e, 'h107e5, 'h103bc, 'h106ed, 'h106f5, 'h1075f, 'h106fd, 'h10705, 'h10760, 'h1070d, 'h10715, 'h10761, 'h1071d, 'h10725, 'h10762, 'h1072d, 'h10735, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h107e5, 'h103bc, 'h10745, 'h10764, 'h1074d, 'h10755, 'h10765, 'h1075d, 'h106e5, 'h10766, 'h107ed, 'h106ed, 'h106f5, 'h10767, 'h106fd, 'h10705, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10769, 'h103bc, 'h1071d, 'h10725, 'h1076a, 'h1072d, 'h10735, 'h1076b, 'h1073d, 'h107ed, 'h10745, 'h1076c, 'h1074d, 'h10755, 'h1076d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1076e, 'h107f5, 'h103bc, 'h106ed, 'h106f5, 'h1076f, 'h106fd, 'h10705, 'h10770, 'h1070d, 'h10715, 'h10771, 'h1071d, 'h10725, 'h10772, 'h1072d, 'h10735, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h107f5, 'h103bc, 'h10745, 'h10774, 'h1074d, 'h10755, 'h10775, 'h1075d, 'h106e5, 'h10776, 'h107fd, 'h106ed, 'h106f5, 'h10777, 'h106fd, 'h10705, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10779, 'h103bc, 'h1071d, 'h10725, 'h1077a, 'h1072d, 'h10735, 'h1077b, 'h1073d, 'h107fd, 'h10745, 'h1077c, 'h1074d, 'h10755, 'h1077d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1077e, 'h10805, 'h103bc, 'h106ed, 'h106f5, 'h1077f, 'h106fd, 'h10705, 'h10780, 'h1070d, 'h10715, 'h10781, 'h1071d, 'h10725, 'h10782, 'h1072d, 'h10735, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10805, 'h103bc, 'h10745, 'h10784, 'h1074d, 'h10755, 'h10785, 'h1075d, 'h106e5, 'h10786, 'h1080d, 'h106ed, 'h106f5, 'h10787, 'h106fd, 'h10705, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10789, 'h103bc, 'h1071d, 'h10725, 'h1078a, 'h1072d, 'h10735, 'h1078b, 'h1073d, 'h1080d, 'h10745, 'h1078c, 'h1074d, 'h10755, 'h1078d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1078e, 'h10815, 'h103bc, 'h106ed, 'h106f5, 'h1078f, 'h106fd, 'h10705, 'h10790, 'h1070d, 'h10715, 'h10791, 'h1071d, 'h10725, 'h10792, 'h1072d, 'h10735, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10815, 'h103bc, 'h10745, 'h10794, 'h1074d, 'h10755, 'h10795, 'h1075d, 'h106e5, 'h10796, 'h1081d, 'h106ed, 'h106f5, 'h10797, 'h106fd, 'h10705, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10799, 'h103bc, 'h1071d, 'h10725, 'h1079a, 'h1072d, 'h10735, 'h1079b, 'h1073d, 'h1081d, 'h10745, 'h1079c, 'h1074d, 'h10755, 'h1079d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1079e, 'h10825, 'h103bc, 'h106ed, 'h106f5, 'h1079f, 'h106fd, 'h10705, 'h107a0, 'h1070d, 'h10715, 'h107a1, 'h1071d, 'h10725, 'h107a2, 'h1072d, 'h10735, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10825, 'h103bc, 'h10745, 'h107a4, 'h1074d, 'h10755, 'h107a5, 'h1075d, 'h106e5, 'h107a6, 'h1082d, 'h106ed, 'h106f5, 'h107a7, 'h106fd, 'h10705, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107a9, 'h103bc, 'h1071d, 'h10725, 'h107aa, 'h1072d, 'h10735, 'h107ab, 'h1073d, 'h1082d, 'h10745, 'h107ac, 'h1074d, 'h10755, 'h107ad, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h107ae, 'h10835, 'h103bc, 'h106ed, 'h106f5, 'h107af, 'h106fd, 'h10705, 'h107b0, 'h1070d, 'h10715, 'h107b1, 'h1071d, 'h10725, 'h107b2, 'h1072d, 'h10735, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10835, 'h103bc, 'h10745, 'h107b4, 'h1074d, 'h10755, 'h107b5, 'h1075d, 'h106e5, 'h107b6, 'h1083d, 'h106ed, 'h106f5, 'h107b7, 'h106fd, 'h10705, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107b9, 'h103bc, 'h1071d, 'h10725, 'h107ba, 'h1072d, 'h10735, 'h107bb, 'h1073d, 'h1083d, 'h10745, 'h107bc, 'h1074d, 'h10755, 'h107bd, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h107be, 'h10845, 'h103bc, 'h106ed, 'h106f5, 'h107bf, 'h106fd, 'h10705, 'h107c0, 'h1070d, 'h10715, 'h107c1, 'h1071d, 'h10725, 'h107c2, 'h1072d, 'h10735, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10845, 'h103bc, 'h10745, 'h107c4, 'h1074d, 'h10755, 'h107c5, 'h1075d, 'h106e5, 'h107c6, 'h1084d, 'h106ed, 'h106f5, 'h107c7, 'h106fd, 'h10705, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107c9, 'h103bc, 'h1071d, 'h10725, 'h107ca, 'h1072d, 'h10735, 'h107cb, 'h1073d, 'h1084d, 'h10745, 'h107cc, 'h1074d, 'h10755, 'h107cd, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h107ce, 'h10855, 'h103bc, 'h106ed, 'h106f5, 'h107cf, 'h106fd, 'h10705, 'h107d0, 'h1070d, 'h10715, 'h107d1, 'h1071d, 'h10725, 'h107d2, 'h1072d, 'h10735, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10855, 'h103bc, 'h10745, 'h107d4, 'h1074d, 'h10755, 'h107d5, 'h1075d, 'h106e5, 'h107d6, 'h1085d, 'h106ed, 'h106f5, 'h107d7, 'h106fd, 'h10705, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107d9, 'h103bc, 'h1071d, 'h10725, 'h107da, 'h1072d, 'h10735, 'h107db, 'h1073d, 'h1085d, 'h10745, 'h107dc, 'h1074d, 'h10755, 'h107dd, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1075e, 'h107e5, 'h103bc, 'h106ed, 'h106f5, 'h1075f, 'h106fd, 'h10705, 'h10760, 'h1070d, 'h10715, 'h10761, 'h1071d, 'h10725, 'h10762, 'h1072d, 'h10735, 'h10763, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h107e5, 'h103bc, 'h10745, 'h10764, 'h1074d, 'h10755, 'h10765, 'h1075d, 'h106e5, 'h10766, 'h107ed, 'h106ed, 'h106f5, 'h10767, 'h106fd, 'h10705, 'h10768, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10769, 'h103bc, 'h1071d, 'h10725, 'h1076a, 'h1072d, 'h10735, 'h1076b, 'h1073d, 'h107ed, 'h10745, 'h1076c, 'h1074d, 'h10755, 'h1076d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1076e, 'h107f5, 'h103bc, 'h106ed, 'h106f5, 'h1076f, 'h106fd, 'h10705, 'h10770, 'h1070d, 'h10715, 'h10771, 'h1071d, 'h10725, 'h10772, 'h1072d, 'h10735, 'h10773, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h107f5, 'h103bc, 'h10745, 'h10774, 'h1074d, 'h10755, 'h10775, 'h1075d, 'h106e5, 'h10776, 'h107fd, 'h106ed, 'h106f5, 'h10777, 'h106fd, 'h10705, 'h10778, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10779, 'h103bc, 'h1071d, 'h10725, 'h1077a, 'h1072d, 'h10735, 'h1077b, 'h1073d, 'h107fd, 'h10745, 'h1077c, 'h1074d, 'h10755, 'h1077d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1077e, 'h10805, 'h103bc, 'h106ed, 'h106f5, 'h1077f, 'h106fd, 'h10705, 'h10780, 'h1070d, 'h10715, 'h10781, 'h1071d, 'h10725, 'h10782, 'h1072d, 'h10735, 'h10783, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10805, 'h103bc, 'h10745, 'h10784, 'h1074d, 'h10755, 'h10785, 'h1075d, 'h106e5, 'h10786, 'h1080d, 'h106ed, 'h106f5, 'h10787, 'h106fd, 'h10705, 'h10788, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10789, 'h103bc, 'h1071d, 'h10725, 'h1078a, 'h1072d, 'h10735, 'h1078b, 'h1073d, 'h1080d, 'h10745, 'h1078c, 'h1074d, 'h10755, 'h1078d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1078e, 'h10815, 'h103bc, 'h106ed, 'h106f5, 'h1078f, 'h106fd, 'h10705, 'h10790, 'h1070d, 'h10715, 'h10791, 'h1071d, 'h10725, 'h10792, 'h1072d, 'h10735, 'h10793, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10815, 'h103bc, 'h10745, 'h10794, 'h1074d, 'h10755, 'h10795, 'h1075d, 'h106e5, 'h10796, 'h1081d, 'h106ed, 'h106f5, 'h10797, 'h106fd, 'h10705, 'h10798, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h10799, 'h103bc, 'h1071d, 'h10725, 'h1079a, 'h1072d, 'h10735, 'h1079b, 'h1073d, 'h1081d, 'h10745, 'h1079c, 'h1074d, 'h10755, 'h1079d, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h1079e, 'h10825, 'h103bc, 'h106ed, 'h106f5, 'h1079f, 'h106fd, 'h10705, 'h107a0, 'h1070d, 'h10715, 'h107a1, 'h1071d, 'h10725, 'h107a2, 'h1072d, 'h10735, 'h107a3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10825, 'h103bc, 'h10745, 'h107a4, 'h1074d, 'h10755, 'h107a5, 'h1075d, 'h106e5, 'h107a6, 'h1082d, 'h106ed, 'h106f5, 'h107a7, 'h106fd, 'h10705, 'h107a8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107a9, 'h103bc, 'h1071d, 'h10725, 'h107aa, 'h1072d, 'h10735, 'h107ab, 'h1073d, 'h1082d, 'h10745, 'h107ac, 'h1074d, 'h10755, 'h107ad, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h107ae, 'h10835, 'h103bc, 'h106ed, 'h106f5, 'h107af, 'h106fd, 'h10705, 'h107b0, 'h1070d, 'h10715, 'h107b1, 'h1071d, 'h10725, 'h107b2, 'h1072d, 'h10735, 'h107b3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10835, 'h103bc, 'h10745, 'h107b4, 'h1074d, 'h10755, 'h107b5, 'h1075d, 'h106e5, 'h107b6, 'h1083d, 'h106ed, 'h106f5, 'h107b7, 'h106fd, 'h10705, 'h107b8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107b9, 'h103bc, 'h1071d, 'h10725, 'h107ba, 'h1072d, 'h10735, 'h107bb, 'h1073d, 'h1083d, 'h10745, 'h107bc, 'h1074d, 'h10755, 'h107bd, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h107be, 'h10845, 'h103bc, 'h106ed, 'h106f5, 'h107bf, 'h106fd, 'h10705, 'h107c0, 'h1070d, 'h10715, 'h107c1, 'h1071d, 'h10725, 'h107c2, 'h1072d, 'h10735, 'h107c3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10845, 'h103bc, 'h10745, 'h107c4, 'h1074d, 'h10755, 'h107c5, 'h1075d, 'h106e5, 'h107c6, 'h1084d, 'h106ed, 'h106f5, 'h107c7, 'h106fd, 'h10705, 'h107c8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107c9, 'h103bc, 'h1071d, 'h10725, 'h107ca, 'h1072d, 'h10735, 'h107cb, 'h1073d, 'h1084d, 'h10745, 'h107cc, 'h1074d, 'h10755, 'h107cd, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h107ce, 'h10855, 'h103bc, 'h106ed, 'h106f5, 'h107cf, 'h106fd, 'h10705, 'h107d0, 'h1070d, 'h10715, 'h107d1, 'h1071d, 'h10725, 'h107d2, 'h1072d, 'h10735, 'h107d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h1073d, 'h10855, 'h103bc, 'h10745, 'h107d4, 'h1074d, 'h10755, 'h107d5, 'h1075d, 'h106e5, 'h107d6, 'h1085d, 'h106ed, 'h106f5, 'h107d7, 'h106fd, 'h10705, 'h107d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h1070d, 'h10715, 'h107d9, 'h103bc, 'h1071d, 'h10725, 'h107da, 'h1072d, 'h10735, 'h107db, 'h1073d, 'h1085d, 'h10745, 'h107dc, 'h1074d, 'h10755, 'h107dd, 'h1075d, 'h21f8e, 'h21f8f, 'h21f8c, 'h21f8b, 'h21f8d, 'h10440, 'h21f8a, 'h10443, 'h10442, 'h1043f, 'h10441, 'h103dc, 'h103dd, 'h21f88, 'h21f89, 'h21f87, 'h103de, 'h103df, 'h103e0, 'h103e1, 'h103e2, 'h103e3, 'h103e4, 'h103e5, 'h103e6, 'h103e7, 'h103e8, 'h103e9, 'h103ea, 'h103eb, 'h103ec, 'h103ed, 'h103ee, 'h103ef, 'h103f0, 'h103f1, 'h103f2, 'h103f3, 'h103f4, 'h103f5, 'h103f6, 'h103f7, 'h103f8, 'h103f9, 'h103fa, 'h103fb, 'h103fc, 'h103fd, 'h103fe, 'h103ff, 'h10400, 'h10401, 'h10402, 'h10403, 'h10404, 'h10405, 'h10406, 'h10407, 'h10408, 'h10409, 'h1040a, 'h1040b, 'h1040c, 'h1040d, 'h1040e, 'h1040f, 'h10410, 'h10411, 'h10412, 'h10413, 'h10414, 'h10415, 'h10416, 'h10417, 'h10418, 'h10419, 'h1041a, 'h1041b, 'h1041c, 'h1041d, 'h1041e, 'h1041f, 'h10420, 'h10421, 'h10422, 'h10423, 'h10424, 'h10425, 'h10426, 'h10427, 'h10428, 'h10429, 'h1042a, 'h1042b, 'h1042c, 'h1042d, 'h1042e, 'h1042f, 'h10430, 'h10431, 'h10432, 'h10433, 'h10434, 'h10435, 'h10436, 'h10437, 'h10438, 'h10439, 'h1043a, 'h1043b, 'h1043c, 'h1043d, 'h1043e, 'h1043f, 'h10442, 'h21f8c, 'h21f8a, 'h21f8b, 'h21f8d, 'h21f8f};;
	
endpackage