

package TESTCASES;
	
	import QSORT_PKG::QSORT_DATA, QSORT_PKG::QSORT_DATA_SIZE, MATRIX_MULTIPLY_16_PKG::MM16_DATA, MATRIX_MULTIPLY_16_PKG::MM16_DATA_SIZE, MATRIX_MULTIPLY_32_PKG::MM32_DATA, MATRIX_MULTIPLY_32_PKG::MM32_DATA_SIZE, LU_PKG::LU_DATA, LU_PKG::LU_DATA_SIZE;
	
	parameter TESTCASE_DATA_SIZE = MM16_DATA_SIZE;
	
	int hit_count = 0, miss_count = 0;
	
	int TESTCASE_DATA [TESTCASE_DATA_SIZE-1:0] = MM16_DATA;
	
endpackage