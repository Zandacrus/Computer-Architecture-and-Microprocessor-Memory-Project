

package QSORT_PKG;
	
	parameter QSORT_DATA_SIZE = 524;
	
	int QSORT_DATA [QSORT_DATA_SIZE-1:0] = {'h21f86, 'h103ad, 'h106a0, 'h21f85, 'h21f71, 'h21f74, 'h1042f, 'h21f6d, 'h21f6e, 'h21f70, 'h103c8, 'h103c7, 'h21f60, 'h21f6b, 'h103ae, 'h21f61, 'h21f6a, 'h10440, 'h10498, 'h21f75, 'h10499, 'h21f76, 'h1049a, 'h10003, 'h10002, 'h21f71, 'h21f74, 'h1042f, 'h21f6d, 'h21f6e, 'h21f70, 'h103c8, 'h103c7, 'h1049b, 'h1049c, 'h21f72, 'h103ae, 'h1049d, 'h1049e, 'h1049f, 'h21f75, 'h104a0, 'h21f76, 'h104a1, 'h104a2, 'h10003, 'h10002, 'h21f74, 'h21f71, 'h1042f, 'h21f6d, 'h21f6e, 'h21f70, 'h103c8, 'h103c7, 'h104a3, 'h104a4, 'h21f73, 'h103ae, 'h104a5, 'h104a6, 'h104a7, 'h21f75, 'h104a8, 'h21f76, 'h104a9, 'h104aa, 'h10003, 'h21f74, 'h10002, 'h21f71, 'h1042f, 'h21f6d, 'h21f6e, 'h21f70, 'h103c8, 'h103c7, 'h104ab, 'h104ac, 'h21f6b, 'h21f6c, 'h21f6a, 'h21f69, 'h21f68, 'h21f67, 'h21f66, 'h21f73, 'h21f72, 'h21f65, 'h21f63, 'h21f62, 'h21f61, 'h21f64, 'h21f71, 'h21f74, 'h21f6d, 'h1042f, 'h21f6e, 'h21f70, 'h103c9, 'h21f6f, 'h21f2c, 'h21f2b, 'h21f2a, 'h21f29, 'h21f6c, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h21f1c, 'h21f27, 'h103ae, 'h21f1d, 'h21f6d, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h10599, 'h21f6c, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f72, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h10599, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f72, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h10599, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f72, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h10599, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f72, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h10599, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f73, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h10599, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f73, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h10599, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f73, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h10599, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f73, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f53, 'h21f6c, 'h1059a, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h1042f, 'h21f6d, 'h21f4d, 'h21f4c, 'h21f43, 'h21f30, 'h21f4b, 'h103c8, 'h103ae, 'h21f6b, 'h103ab, 'h21f51, 'h21f50, 'h1008a, 'h21f70, 'h21f4f, 'h21f3c, 'h21f6c, 'h10070, 'h1006f, 'h1006e, 'h21f53, 'h21f6d, 'h1059a, 'h21f6e, 'h103c9, 'h21f2c, 'h21f29, 'h21f2a, 'h21f2b, 'h21f6f, 'h21f74, 'h21f71, 'h21f84, 'h1042c, 'h21f82, 'h21f80, 'h21f81, 'h21f7f, 'h1042f, 'h1042e, 'h1042b, 'h1042d, 'h103c8, 'h21f7d, 'h21f7e, 'h21f7c, 'h103c9, 'h21f7b, 'h21f7a, 'h103ae, 'h1043a, 'h103ca, 'h103cb, 'h103cc, 'h103cd, 'h103ce, 'h103cf, 'h103d0, 'h103d1, 'h103d2, 'h103d3, 'h103d4, 'h103d5, 'h103d6, 'h103d7, 'h103d8, 'h103d9, 'h103da, 'h103db, 'h103dc, 'h103dd, 'h103de, 'h103df, 'h103e0, 'h103e1, 'h103e2, 'h103e3, 'h103e4, 'h103e5, 'h103e6, 'h103e7, 'h103e8, 'h103e9, 'h103ea, 'h103eb, 'h103ec, 'h103ed, 'h103ee, 'h103ef, 'h103f0, 'h103f1, 'h103f2, 'h103f3, 'h103f4, 'h103f5, 'h103f6, 'h103f7, 'h103f8, 'h103f9, 'h103fa, 'h103fb, 'h103fc, 'h103fd, 'h103fe, 'h103ff, 'h10400, 'h10401, 'h10402, 'h10403, 'h10404, 'h10405, 'h10406, 'h10407, 'h10408, 'h10409, 'h1040a, 'h1040b, 'h1040c, 'h1040d, 'h1040e, 'h1040f, 'h10410, 'h10411, 'h10412, 'h10413, 'h10414, 'h10415, 'h10416, 'h10417, 'h10418, 'h10419, 'h1041a, 'h1041b, 'h1041c, 'h1041d, 'h1041e, 'h1041f, 'h10420, 'h10421, 'h10422, 'h10423, 'h10424, 'h10425, 'h10426, 'h10427, 'h10428, 'h10429, 'h1042a, 'h1042b, 'h1042e, 'h21f81, 'h21f7f, 'h21f80, 'h21f82, 'h21f84};
	
endpackage