

package MATRIX_MULTIPLY_32_PKG_5;
	
	import MATRIX_MULTIPLY_32_PKG_4::DATA4;
	
	parameter SIZE = 8500;
	
	int DATA0 [SIZE-1:0] = {'h10775, 'h10785, 'h109d3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10795, 'h10bd5, 'h107a5, 'h109d4, 'h107b5, 'h107c5, 'h109d5, 'h107d5, 'h107e5, 'h109d6, 'h107f5, 'h10805, 'h109d7, 'h10815, 'h103bc, 'h10825, 'h109d8, 'h10835, 'h21f8e, 'h21f8f, 'h21f8d, 'h10845, 'h109d9, 'h10bd5, 'h10855, 'h10865, 'h109da, 'h10875, 'h10885, 'h109db, 'h10895, 'h108a5, 'h109dc, 'h108b5, 'h108c5, 'h109dd, 'h103bc, 'h108d5, 'h106e5, 'h109de, 'h10be5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f5, 'h10705, 'h109df, 'h10715, 'h10725, 'h109e0, 'h10735, 'h10745, 'h109e1, 'h10755, 'h10765, 'h109e2, 'h10775, 'h103bc, 'h10785, 'h109e3, 'h10795, 'h10be5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a5, 'h109e4, 'h107b5, 'h107c5, 'h109e5, 'h107d5, 'h107e5, 'h109e6, 'h107f5, 'h10805, 'h109e7, 'h10815, 'h10825, 'h109e8, 'h103bc, 'h10835, 'h10845, 'h109e9, 'h10be5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10855, 'h10865, 'h109ea, 'h10875, 'h10885, 'h109eb, 'h10895, 'h108a5, 'h109ec, 'h108b5, 'h108c5, 'h109ed, 'h108d5, 'h103bc, 'h106e5, 'h109ee, 'h10bf5, 'h106f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10705, 'h109ef, 'h10715, 'h10725, 'h109f0, 'h10735, 'h10745, 'h109f1, 'h10755, 'h10765, 'h109f2, 'h10775, 'h10785, 'h109f3, 'h103bc, 'h10795, 'h10bf5, 'h107a5, 'h109f4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b5, 'h107c5, 'h109f5, 'h107d5, 'h107e5, 'h109f6, 'h107f5, 'h10805, 'h109f7, 'h10815, 'h10825, 'h109f8, 'h10835, 'h103bc, 'h10845, 'h109f9, 'h10bf5, 'h10855, 'h21f8e, 'h21f8f, 'h21f8d, 'h10865, 'h109fa, 'h10875, 'h10885, 'h109fb, 'h10895, 'h108a5, 'h109fc, 'h108b5, 'h108c5, 'h109fd, 'h108d5, 'h106e5, 'h109fe, 'h10c05, 'h103bc, 'h106f5, 'h10705, 'h109ff, 'h21f8e, 'h21f8f, 'h21f8d, 'h10715, 'h10725, 'h10a00, 'h10735, 'h10745, 'h10a01, 'h10755, 'h10765, 'h10a02, 'h10775, 'h10785, 'h10a03, 'h10795, 'h10c05, 'h103bc, 'h107a5, 'h10a04, 'h107b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c5, 'h10a05, 'h107d5, 'h107e5, 'h10a06, 'h107f5, 'h10805, 'h10a07, 'h10815, 'h10825, 'h10a08, 'h10835, 'h10845, 'h10a09, 'h10c05, 'h103bc, 'h10855, 'h10865, 'h10a0a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10875, 'h10885, 'h10a0b, 'h10895, 'h108a5, 'h10a0c, 'h108b5, 'h108c5, 'h10a0d, 'h108d5, 'h106e5, 'h10a0e, 'h10c15, 'h106f5, 'h103bc, 'h10705, 'h10a0f, 'h10715, 'h21f8e, 'h21f8f, 'h21f8d, 'h10725, 'h10a10, 'h10735, 'h10745, 'h10a11, 'h10755, 'h10765, 'h10a12, 'h10775, 'h10785, 'h10a13, 'h10795, 'h10c15, 'h107a5, 'h10a14, 'h103bc, 'h107b5, 'h107c5, 'h10a15, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d5, 'h107e5, 'h10a16, 'h107f5, 'h10805, 'h10a17, 'h10815, 'h10825, 'h10a18, 'h10835, 'h10845, 'h10a19, 'h10c15, 'h10855, 'h103bc, 'h10865, 'h10a1a, 'h10875, 'h21f8e, 'h21f8f, 'h21f8d, 'h10885, 'h10a1b, 'h10895, 'h108a5, 'h10a1c, 'h108b5, 'h108c5, 'h10a1d, 'h108d5, 'h106e5, 'h10a1e, 'h10c25, 'h106f5, 'h10705, 'h10a1f, 'h103bc, 'h10715, 'h10725, 'h10a20, 'h21f8e, 'h21f8f, 'h21f8d, 'h10735, 'h10745, 'h10a21, 'h10755, 'h10765, 'h10a22, 'h10775, 'h10785, 'h10a23, 'h10795, 'h10c25, 'h107a5, 'h10a24, 'h107b5, 'h103bc, 'h107c5, 'h10a25, 'h107d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e5, 'h10a26, 'h107f5, 'h10805, 'h10a27, 'h10815, 'h10825, 'h10a28, 'h10835, 'h10845, 'h10a29, 'h10c25, 'h10855, 'h10865, 'h10a2a, 'h103bc, 'h10875, 'h10885, 'h10a2b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10895, 'h108a5, 'h10a2c, 'h108b5, 'h108c5, 'h10a2d, 'h108d5, 'h106e5, 'h10a2e, 'h10c35, 'h106f5, 'h10705, 'h10a2f, 'h10715, 'h103bc, 'h10725, 'h10a30, 'h10735, 'h21f8e, 'h21f8f, 'h21f8d, 'h10745, 'h10a31, 'h10755, 'h10765, 'h10a32, 'h10775, 'h10785, 'h10a33, 'h10795, 'h10c35, 'h107a5, 'h10a34, 'h107b5, 'h107c5, 'h10a35, 'h103bc, 'h107d5, 'h107e5, 'h10a36, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f5, 'h10805, 'h10a37, 'h10815, 'h10825, 'h10a38, 'h10835, 'h10845, 'h10a39, 'h10c35, 'h10855, 'h10865, 'h10a3a, 'h10875, 'h103bc, 'h10885, 'h10a3b, 'h10895, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a5, 'h10a3c, 'h108b5, 'h108c5, 'h10a3d, 'h108d5, 'h106e5, 'h10a3e, 'h10c45, 'h106f5, 'h10705, 'h10a3f, 'h10715, 'h10725, 'h10a40, 'h103bc, 'h10735, 'h10745, 'h10a41, 'h21f8e, 'h21f8f, 'h21f8d, 'h10755, 'h10765, 'h10a42, 'h10775, 'h10785, 'h10a43, 'h10795, 'h10c45, 'h107a5, 'h10a44, 'h107b5, 'h107c5, 'h10a45, 'h107d5, 'h103bc, 'h107e5, 'h10a46, 'h107f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10805, 'h10a47, 'h10815, 'h10825, 'h10a48, 'h10835, 'h10845, 'h10a49, 'h10c45, 'h10855, 'h10865, 'h10a4a, 'h10875, 'h10885, 'h10a4b, 'h103bc, 'h10895, 'h108a5, 'h10a4c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b5, 'h108c5, 'h10a4d, 'h108d5, 'h106e5, 'h10a4e, 'h10c55, 'h106f5, 'h10705, 'h10a4f, 'h10715, 'h10725, 'h10a50, 'h10735, 'h103bc, 'h10745, 'h10a51, 'h10755, 'h21f8e, 'h21f8f, 'h21f8d, 'h10765, 'h10a52, 'h10775, 'h10785, 'h10a53, 'h10795, 'h10c55, 'h107a5, 'h10a54, 'h107b5, 'h107c5, 'h10a55, 'h107d5, 'h107e5, 'h10a56, 'h103bc, 'h107f5, 'h10805, 'h10a57, 'h21f8e, 'h21f8f, 'h21f8d, 'h10815, 'h10825, 'h10a58, 'h10835, 'h10845, 'h10a59, 'h10c55, 'h10855, 'h10865, 'h10a5a, 'h10875, 'h10885, 'h10a5b, 'h10895, 'h103bc, 'h108a5, 'h10a5c, 'h108b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c5, 'h10a5d, 'h108d5, 'h106e5, 'h10a5e, 'h10c65, 'h106f5, 'h10705, 'h10a5f, 'h10715, 'h10725, 'h10a60, 'h10735, 'h10745, 'h10a61, 'h103bc, 'h10755, 'h10765, 'h10a62, 'h21f8e, 'h21f8f, 'h21f8d, 'h10775, 'h10785, 'h10a63, 'h10795, 'h10c65, 'h107a5, 'h10a64, 'h107b5, 'h107c5, 'h10a65, 'h107d5, 'h107e5, 'h10a66, 'h107f5, 'h103bc, 'h10805, 'h10a67, 'h10815, 'h21f8e, 'h21f8f, 'h21f8d, 'h10825, 'h10a68, 'h10835, 'h10845, 'h10a69, 'h10c65, 'h10855, 'h10865, 'h10a6a, 'h10875, 'h10885, 'h10a6b, 'h10895, 'h108a5, 'h10a6c, 'h103bc, 'h108b5, 'h108c5, 'h10a6d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d5, 'h106e5, 'h10a6e, 'h10c75, 'h106f5, 'h10705, 'h10a6f, 'h10715, 'h10725, 'h10a70, 'h10735, 'h10745, 'h10a71, 'h10755, 'h103bc, 'h10765, 'h10a72, 'h10775, 'h21f8e, 'h21f8f, 'h21f8d, 'h10785, 'h10a73, 'h10795, 'h10c75, 'h107a5, 'h10a74, 'h107b5, 'h107c5, 'h10a75, 'h107d5, 'h107e5, 'h10a76, 'h107f5, 'h10805, 'h10a77, 'h103bc, 'h10815, 'h10825, 'h10a78, 'h21f8e, 'h21f8f, 'h21f8d, 'h10835, 'h10845, 'h10a79, 'h10c75, 'h10855, 'h10865, 'h10a7a, 'h10875, 'h10885, 'h10a7b, 'h10895, 'h108a5, 'h10a7c, 'h108b5, 'h103bc, 'h108c5, 'h10a7d, 'h108d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e5, 'h10a7e, 'h10c85, 'h106f5, 'h10705, 'h10a7f, 'h10715, 'h10725, 'h10a80, 'h10735, 'h10745, 'h10a81, 'h10755, 'h10765, 'h10a82, 'h103bc, 'h10775, 'h10785, 'h10a83, 'h21f8e, 'h21f8f, 'h21f8d, 'h10795, 'h10c85, 'h107a5, 'h10a84, 'h107b5, 'h107c5, 'h10a85, 'h107d5, 'h107e5, 'h10a86, 'h107f5, 'h10805, 'h10a87, 'h10815, 'h103bc, 'h10825, 'h10a88, 'h10835, 'h21f8e, 'h21f8f, 'h21f8d, 'h10845, 'h10a89, 'h10c85, 'h10855, 'h10865, 'h10a8a, 'h10875, 'h10885, 'h10a8b, 'h10895, 'h108a5, 'h10a8c, 'h108b5, 'h108c5, 'h10a8d, 'h103bc, 'h108d5, 'h106e5, 'h10a8e, 'h10c95, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f5, 'h10705, 'h10a8f, 'h10715, 'h10725, 'h10a90, 'h10735, 'h10745, 'h10a91, 'h10755, 'h10765, 'h10a92, 'h10775, 'h103bc, 'h10785, 'h10a93, 'h10795, 'h10c95, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a5, 'h10a94, 'h107b5, 'h107c5, 'h10a95, 'h107d5, 'h107e5, 'h10a96, 'h107f5, 'h10805, 'h10a97, 'h10815, 'h10825, 'h10a98, 'h103bc, 'h10835, 'h10845, 'h10a99, 'h10c95, 'h21f8e, 'h21f8f, 'h21f8d, 'h10855, 'h10865, 'h10a9a, 'h10875, 'h10885, 'h10a9b, 'h10895, 'h108a5, 'h10a9c, 'h108b5, 'h108c5, 'h10a9d, 'h108d5, 'h103bc, 'h106e5, 'h10a9e, 'h10ca5, 'h106f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h10705, 'h10a9f, 'h10715, 'h10725, 'h10aa0, 'h10735, 'h10745, 'h10aa1, 'h10755, 'h10765, 'h10aa2, 'h10775, 'h10785, 'h10aa3, 'h103bc, 'h10795, 'h10ca5, 'h107a5, 'h10aa4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b5, 'h107c5, 'h10aa5, 'h107d5, 'h107e5, 'h10aa6, 'h107f5, 'h10805, 'h10aa7, 'h10815, 'h10825, 'h10aa8, 'h10835, 'h103bc, 'h10845, 'h10aa9, 'h10ca5, 'h10855, 'h21f8e, 'h21f8f, 'h21f8d, 'h10865, 'h10aaa, 'h10875, 'h10885, 'h10aab, 'h10895, 'h108a5, 'h10aac, 'h108b5, 'h108c5, 'h10aad, 'h108d5, 'h106e5, 'h10aae, 'h10cb5, 'h103bc, 'h106f5, 'h10705, 'h10aaf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10715, 'h10725, 'h10ab0, 'h10735, 'h10745, 'h10ab1, 'h10755, 'h10765, 'h10ab2, 'h10775, 'h10785, 'h10ab3, 'h10795, 'h10cb5, 'h103bc, 'h107a5, 'h10ab4, 'h107b5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c5, 'h10ab5, 'h107d5, 'h107e5, 'h10ab6, 'h107f5, 'h10805, 'h10ab7, 'h10815, 'h10825, 'h10ab8, 'h10835, 'h10845, 'h10ab9, 'h10cb5, 'h103bc, 'h10855, 'h10865, 'h10aba, 'h21f8e, 'h21f8f, 'h21f8d, 'h10875, 'h10885, 'h10abb, 'h10895, 'h108a5, 'h10abc, 'h108b5, 'h108c5, 'h10abd, 'h108d5, 'h106e5, 'h10abe, 'h10cc5, 'h106f5, 'h103bc, 'h10705, 'h10abf, 'h10715, 'h21f8e, 'h21f8f, 'h21f8d, 'h10725, 'h10ac0, 'h10735, 'h10745, 'h10ac1, 'h10755, 'h10765, 'h10ac2, 'h10775, 'h10785, 'h10ac3, 'h10795, 'h10cc5, 'h107a5, 'h10ac4, 'h103bc, 'h107b5, 'h107c5, 'h10ac5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d5, 'h107e5, 'h10ac6, 'h107f5, 'h10805, 'h10ac7, 'h10815, 'h10825, 'h10ac8, 'h10835, 'h10845, 'h10ac9, 'h10cc5, 'h10855, 'h103bc, 'h10865, 'h10aca, 'h10875, 'h21f8e, 'h21f8f, 'h21f8d, 'h10885, 'h10acb, 'h10895, 'h108a5, 'h10acc, 'h108b5, 'h108c5, 'h10acd, 'h108d5, 'h106e5, 'h10ace, 'h10cd5, 'h106f5, 'h10705, 'h10acf, 'h103bc, 'h10715, 'h10725, 'h10ad0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10735, 'h10745, 'h10ad1, 'h10755, 'h10765, 'h10ad2, 'h10775, 'h10785, 'h10ad3, 'h10795, 'h10cd5, 'h107a5, 'h10ad4, 'h107b5, 'h103bc, 'h107c5, 'h10ad5, 'h107d5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e5, 'h10ad6, 'h107f5, 'h10805, 'h10ad7, 'h10815, 'h10825, 'h10ad8, 'h10835, 'h10845, 'h10ad9, 'h10cd5, 'h10855, 'h10865, 'h10ada, 'h103bc, 'h10875, 'h10885, 'h10adb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10895, 'h108a5, 'h10adc, 'h108b5, 'h108c5, 'h10add, 'h108d5, 'h106e6, 'h108de, 'h10ae6, 'h106f6, 'h10706, 'h108df, 'h10716, 'h103bc, 'h10726, 'h108e0, 'h10736, 'h21f8e, 'h21f8f, 'h21f8d, 'h10746, 'h108e1, 'h10756, 'h10766, 'h108e2, 'h10776, 'h10786, 'h108e3, 'h10796, 'h10ae6, 'h107a6, 'h108e4, 'h107b6, 'h107c6, 'h108e5, 'h103bc, 'h107d6, 'h107e6, 'h108e6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f6, 'h10806, 'h108e7, 'h10816, 'h10826, 'h108e8, 'h10836, 'h10846, 'h108e9, 'h10ae6, 'h10856, 'h10866, 'h108ea, 'h10876, 'h103bc, 'h10886, 'h108eb, 'h10896, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a6, 'h108ec, 'h108b6, 'h108c6, 'h108ed, 'h108d6, 'h106e6, 'h108ee, 'h10af6, 'h106f6, 'h10706, 'h108ef, 'h10716, 'h10726, 'h108f0, 'h103bc, 'h10736, 'h10746, 'h108f1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10756, 'h10766, 'h108f2, 'h10776, 'h10786, 'h108f3, 'h10796, 'h10af6, 'h107a6, 'h108f4, 'h107b6, 'h107c6, 'h108f5, 'h107d6, 'h103bc, 'h107e6, 'h108f6, 'h107f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10806, 'h108f7, 'h10816, 'h10826, 'h108f8, 'h10836, 'h10846, 'h108f9, 'h10af6, 'h10856, 'h10866, 'h108fa, 'h10876, 'h10886, 'h108fb, 'h103bc, 'h10896, 'h108a6, 'h108fc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b6, 'h108c6, 'h108fd, 'h108d6, 'h106e6, 'h108fe, 'h10b06, 'h106f6, 'h10706, 'h108ff, 'h10716, 'h10726, 'h10900, 'h10736, 'h103bc, 'h10746, 'h10901, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h10766, 'h10902, 'h10776, 'h10786, 'h10903, 'h10796, 'h10b06, 'h107a6, 'h10904, 'h107b6, 'h107c6, 'h10905, 'h107d6, 'h107e6, 'h10906, 'h103bc, 'h107f6, 'h10806, 'h10907, 'h21f8e, 'h21f8f, 'h21f8d, 'h10816, 'h10826, 'h10908, 'h10836, 'h10846, 'h10909, 'h10b06, 'h10856, 'h10866, 'h1090a, 'h10876, 'h10886, 'h1090b, 'h10896, 'h103bc, 'h108a6, 'h1090c, 'h108b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c6, 'h1090d, 'h108d6, 'h106e6, 'h1090e, 'h10b16, 'h106f6, 'h10706, 'h1090f, 'h10716, 'h10726, 'h10910, 'h10736, 'h10746, 'h10911, 'h103bc, 'h10756, 'h10766, 'h10912, 'h21f8e, 'h21f8f, 'h21f8d, 'h10776, 'h10786, 'h10913, 'h10796, 'h10b16, 'h107a6, 'h10914, 'h107b6, 'h107c6, 'h10915, 'h107d6, 'h107e6, 'h10916, 'h107f6, 'h103bc, 'h10806, 'h10917, 'h10816, 'h21f8e, 'h21f8f, 'h21f8d, 'h10826, 'h10918, 'h10836, 'h10846, 'h10919, 'h10b16, 'h10856, 'h10866, 'h1091a, 'h10876, 'h10886, 'h1091b, 'h10896, 'h108a6, 'h1091c, 'h103bc, 'h108b6, 'h108c6, 'h1091d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d6, 'h106e6, 'h1091e, 'h10b26, 'h106f6, 'h10706, 'h1091f, 'h10716, 'h10726, 'h10920, 'h10736, 'h10746, 'h10921, 'h10756, 'h103bc, 'h10766, 'h10922, 'h10776, 'h21f8e, 'h21f8f, 'h21f8d, 'h10786, 'h10923, 'h10796, 'h10b26, 'h107a6, 'h10924, 'h107b6, 'h107c6, 'h10925, 'h107d6, 'h107e6, 'h10926, 'h107f6, 'h10806, 'h10927, 'h103bc, 'h10816, 'h10826, 'h10928, 'h21f8e, 'h21f8f, 'h21f8d, 'h10836, 'h10846, 'h10929, 'h10b26, 'h10856, 'h10866, 'h1092a, 'h10876, 'h10886, 'h1092b, 'h10896, 'h108a6, 'h1092c, 'h108b6, 'h103bc, 'h108c6, 'h1092d, 'h108d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e6, 'h1092e, 'h10b36, 'h106f6, 'h10706, 'h1092f, 'h10716, 'h10726, 'h10930, 'h10736, 'h10746, 'h10931, 'h10756, 'h10766, 'h10932, 'h103bc, 'h10776, 'h10786, 'h10933, 'h21f8e, 'h21f8f, 'h21f8d, 'h10796, 'h10b36, 'h107a6, 'h10934, 'h107b6, 'h107c6, 'h10935, 'h107d6, 'h107e6, 'h10936, 'h107f6, 'h10806, 'h10937, 'h10816, 'h103bc, 'h10826, 'h10938, 'h10836, 'h21f8e, 'h21f8f, 'h21f8d, 'h10846, 'h10939, 'h10b36, 'h10856, 'h10866, 'h1093a, 'h10876, 'h10886, 'h1093b, 'h10896, 'h108a6, 'h1093c, 'h108b6, 'h108c6, 'h1093d, 'h103bc, 'h108d6, 'h106e6, 'h1093e, 'h10b46, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f6, 'h10706, 'h1093f, 'h10716, 'h10726, 'h10940, 'h10736, 'h10746, 'h10941, 'h10756, 'h10766, 'h10942, 'h10776, 'h103bc, 'h10786, 'h10943, 'h10796, 'h10b46, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a6, 'h10944, 'h107b6, 'h107c6, 'h10945, 'h107d6, 'h107e6, 'h10946, 'h107f6, 'h10806, 'h10947, 'h10816, 'h10826, 'h10948, 'h103bc, 'h10836, 'h10846, 'h10949, 'h10b46, 'h21f8e, 'h21f8f, 'h21f8d, 'h10856, 'h10866, 'h1094a, 'h10876, 'h10886, 'h1094b, 'h10896, 'h108a6, 'h1094c, 'h108b6, 'h108c6, 'h1094d, 'h108d6, 'h103bc, 'h106e6, 'h1094e, 'h10b56, 'h106f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1094f, 'h10716, 'h10726, 'h10950, 'h10736, 'h10746, 'h10951, 'h10756, 'h10766, 'h10952, 'h10776, 'h10786, 'h10953, 'h103bc, 'h10796, 'h10b56, 'h107a6, 'h10954, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b6, 'h107c6, 'h10955, 'h107d6, 'h107e6, 'h10956, 'h107f6, 'h10806, 'h10957, 'h10816, 'h10826, 'h10958, 'h10836, 'h103bc, 'h10846, 'h10959, 'h10b56, 'h10856, 'h21f8e, 'h21f8f, 'h21f8d, 'h10866, 'h1095a, 'h10876, 'h10886, 'h1095b, 'h10896, 'h108a6, 'h1095c, 'h108b6, 'h108c6, 'h1095d, 'h108d6, 'h106e6, 'h1095e, 'h10b66, 'h103bc, 'h106f6, 'h10706, 'h1095f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10716, 'h10726, 'h10960, 'h10736, 'h10746, 'h10961, 'h10756, 'h10766, 'h10962, 'h10776, 'h10786, 'h10963, 'h10796, 'h10b66, 'h103bc, 'h107a6, 'h10964, 'h107b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c6, 'h10965, 'h107d6, 'h107e6, 'h10966, 'h107f6, 'h10806, 'h10967, 'h10816, 'h10826, 'h10968, 'h10836, 'h10846, 'h10969, 'h10b66, 'h103bc, 'h10856, 'h10866, 'h1096a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10876, 'h10886, 'h1096b, 'h10896, 'h108a6, 'h1096c, 'h108b6, 'h108c6, 'h1096d, 'h108d6, 'h106e6, 'h1096e, 'h10b76, 'h106f6, 'h103bc, 'h10706, 'h1096f, 'h10716, 'h21f8e, 'h21f8f, 'h21f8d, 'h10726, 'h10970, 'h10736, 'h10746, 'h10971, 'h10756, 'h10766, 'h10972, 'h10776, 'h10786, 'h10973, 'h10796, 'h10b76, 'h107a6, 'h10974, 'h103bc, 'h107b6, 'h107c6, 'h10975, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d6, 'h107e6, 'h10976, 'h107f6, 'h10806, 'h10977, 'h10816, 'h10826, 'h10978, 'h10836, 'h10846, 'h10979, 'h10b76, 'h10856, 'h103bc, 'h10866, 'h1097a, 'h10876, 'h21f8e, 'h21f8f, 'h21f8d, 'h10886, 'h1097b, 'h10896, 'h108a6, 'h1097c, 'h108b6, 'h108c6, 'h1097d, 'h108d6, 'h106e6, 'h1097e, 'h10b86, 'h106f6, 'h10706, 'h1097f, 'h103bc, 'h10716, 'h10726, 'h10980, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h10746, 'h10981, 'h10756, 'h10766, 'h10982, 'h10776, 'h10786, 'h10983, 'h10796, 'h10b86, 'h107a6, 'h10984, 'h107b6, 'h103bc, 'h107c6, 'h10985, 'h107d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e6, 'h10986, 'h107f6, 'h10806, 'h10987, 'h10816, 'h10826, 'h10988, 'h10836, 'h10846, 'h10989, 'h10b86, 'h10856, 'h10866, 'h1098a, 'h103bc, 'h10876, 'h10886, 'h1098b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10896, 'h108a6, 'h1098c, 'h108b6, 'h108c6, 'h1098d, 'h108d6, 'h106e6, 'h1098e, 'h10b96, 'h106f6, 'h10706, 'h1098f, 'h10716, 'h103bc, 'h10726, 'h10990, 'h10736, 'h21f8e, 'h21f8f, 'h21f8d, 'h10746, 'h10991, 'h10756, 'h10766, 'h10992, 'h10776, 'h10786, 'h10993, 'h10796, 'h10b96, 'h107a6, 'h10994, 'h107b6, 'h107c6, 'h10995, 'h103bc, 'h107d6, 'h107e6, 'h10996, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f6, 'h10806, 'h10997, 'h10816, 'h10826, 'h10998, 'h10836, 'h10846, 'h10999, 'h10b96, 'h10856, 'h10866, 'h1099a, 'h10876, 'h103bc, 'h10886, 'h1099b, 'h10896, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a6, 'h1099c, 'h108b6, 'h108c6, 'h1099d, 'h108d6, 'h106e6, 'h1099e, 'h10ba6, 'h106f6, 'h10706, 'h1099f, 'h10716, 'h10726, 'h109a0, 'h103bc, 'h10736, 'h10746, 'h109a1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10756, 'h10766, 'h109a2, 'h10776, 'h10786, 'h109a3, 'h10796, 'h10ba6, 'h107a6, 'h109a4, 'h107b6, 'h107c6, 'h109a5, 'h107d6, 'h103bc, 'h107e6, 'h109a6, 'h107f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10806, 'h109a7, 'h10816, 'h10826, 'h109a8, 'h10836, 'h10846, 'h109a9, 'h10ba6, 'h10856, 'h10866, 'h109aa, 'h10876, 'h10886, 'h109ab, 'h103bc, 'h10896, 'h108a6, 'h109ac, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b6, 'h108c6, 'h109ad, 'h108d6, 'h106e6, 'h109ae, 'h10bb6, 'h106f6, 'h10706, 'h109af, 'h10716, 'h10726, 'h109b0, 'h10736, 'h103bc, 'h10746, 'h109b1, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h10766, 'h109b2, 'h10776, 'h10786, 'h109b3, 'h10796, 'h10bb6, 'h107a6, 'h109b4, 'h107b6, 'h107c6, 'h109b5, 'h107d6, 'h107e6, 'h109b6, 'h103bc, 'h107f6, 'h10806, 'h109b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10816, 'h10826, 'h109b8, 'h10836, 'h10846, 'h109b9, 'h10bb6, 'h10856, 'h10866, 'h109ba, 'h10876, 'h10886, 'h109bb, 'h10896, 'h103bc, 'h108a6, 'h109bc, 'h108b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c6, 'h109bd, 'h108d6, 'h106e6, 'h109be, 'h10bc6, 'h106f6, 'h10706, 'h109bf, 'h10716, 'h10726, 'h109c0, 'h10736, 'h10746, 'h109c1, 'h103bc, 'h10756, 'h10766, 'h109c2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10776, 'h10786, 'h109c3, 'h10796, 'h10bc6, 'h107a6, 'h109c4, 'h107b6, 'h107c6, 'h109c5, 'h107d6, 'h107e6, 'h109c6, 'h107f6, 'h103bc, 'h10806, 'h109c7, 'h10816, 'h21f8e, 'h21f8f, 'h21f8d, 'h10826, 'h109c8, 'h10836, 'h10846, 'h109c9, 'h10bc6, 'h10856, 'h10866, 'h109ca, 'h10876, 'h10886, 'h109cb, 'h10896, 'h108a6, 'h109cc, 'h103bc, 'h108b6, 'h108c6, 'h109cd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d6, 'h106e6, 'h109ce, 'h10bd6, 'h106f6, 'h10706, 'h109cf, 'h10716, 'h10726, 'h109d0, 'h10736, 'h10746, 'h109d1, 'h10756, 'h103bc, 'h10766, 'h109d2, 'h10776, 'h21f8e, 'h21f8f, 'h21f8d, 'h10786, 'h109d3, 'h10796, 'h10bd6, 'h107a6, 'h109d4, 'h107b6, 'h107c6, 'h109d5, 'h107d6, 'h107e6, 'h109d6, 'h107f6, 'h10806, 'h109d7, 'h103bc, 'h10816, 'h10826, 'h109d8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10836, 'h10846, 'h109d9, 'h10bd6, 'h10856, 'h10866, 'h109da, 'h10876, 'h10886, 'h109db, 'h10896, 'h108a6, 'h109dc, 'h108b6, 'h103bc, 'h108c6, 'h109dd, 'h108d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e6, 'h109de, 'h10be6, 'h106f6, 'h10706, 'h109df, 'h10716, 'h10726, 'h109e0, 'h10736, 'h10746, 'h109e1, 'h10756, 'h10766, 'h109e2, 'h103bc, 'h10776, 'h10786, 'h109e3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10796, 'h10be6, 'h107a6, 'h109e4, 'h107b6, 'h107c6, 'h109e5, 'h107d6, 'h107e6, 'h109e6, 'h107f6, 'h10806, 'h109e7, 'h10816, 'h103bc, 'h10826, 'h109e8, 'h10836, 'h21f8e, 'h21f8f, 'h21f8d, 'h10846, 'h109e9, 'h10be6, 'h10856, 'h10866, 'h109ea, 'h10876, 'h10886, 'h109eb, 'h10896, 'h108a6, 'h109ec, 'h108b6, 'h108c6, 'h109ed, 'h103bc, 'h108d6, 'h106e6, 'h109ee, 'h10bf6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f6, 'h10706, 'h109ef, 'h10716, 'h10726, 'h109f0, 'h10736, 'h10746, 'h109f1, 'h10756, 'h10766, 'h109f2, 'h10776, 'h103bc, 'h10786, 'h109f3, 'h10796, 'h10bf6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a6, 'h109f4, 'h107b6, 'h107c6, 'h109f5, 'h107d6, 'h107e6, 'h109f6, 'h107f6, 'h10806, 'h109f7, 'h10816, 'h10826, 'h109f8, 'h103bc, 'h10836, 'h10846, 'h109f9, 'h10bf6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10856, 'h10866, 'h109fa, 'h10876, 'h10886, 'h109fb, 'h10896, 'h108a6, 'h109fc, 'h108b6, 'h108c6, 'h109fd, 'h108d6, 'h103bc, 'h106e6, 'h109fe, 'h10c06, 'h106f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h109ff, 'h10716, 'h10726, 'h10a00, 'h10736, 'h10746, 'h10a01, 'h10756, 'h10766, 'h10a02, 'h10776, 'h10786, 'h10a03, 'h103bc, 'h10796, 'h10c06, 'h107a6, 'h10a04, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b6, 'h107c6, 'h10a05, 'h107d6, 'h107e6, 'h10a06, 'h107f6, 'h10806, 'h10a07, 'h10816, 'h10826, 'h10a08, 'h10836, 'h103bc, 'h10846, 'h10a09, 'h10c06, 'h10856, 'h21f8e, 'h21f8f, 'h21f8d, 'h10866, 'h10a0a, 'h10876, 'h10886, 'h10a0b, 'h10896, 'h108a6, 'h10a0c, 'h108b6, 'h108c6, 'h10a0d, 'h108d6, 'h106e6, 'h10a0e, 'h10c16, 'h103bc, 'h106f6, 'h10706, 'h10a0f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10716, 'h10726, 'h10a10, 'h10736, 'h10746, 'h10a11, 'h10756, 'h10766, 'h10a12, 'h10776, 'h10786, 'h10a13, 'h10796, 'h10c16, 'h103bc, 'h107a6, 'h10a14, 'h107b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c6, 'h10a15, 'h107d6, 'h107e6, 'h10a16, 'h107f6, 'h10806, 'h10a17, 'h10816, 'h10826, 'h10a18, 'h10836, 'h10846, 'h10a19, 'h10c16, 'h103bc, 'h10856, 'h10866, 'h10a1a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10876, 'h10886, 'h10a1b, 'h10896, 'h108a6, 'h10a1c, 'h108b6, 'h108c6, 'h10a1d, 'h108d6, 'h106e6, 'h10a1e, 'h10c26, 'h106f6, 'h103bc, 'h10706, 'h10a1f, 'h10716, 'h21f8e, 'h21f8f, 'h21f8d, 'h10726, 'h10a20, 'h10736, 'h10746, 'h10a21, 'h10756, 'h10766, 'h10a22, 'h10776, 'h10786, 'h10a23, 'h10796, 'h10c26, 'h107a6, 'h10a24, 'h103bc, 'h107b6, 'h107c6, 'h10a25, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d6, 'h107e6, 'h10a26, 'h107f6, 'h10806, 'h10a27, 'h10816, 'h10826, 'h10a28, 'h10836, 'h10846, 'h10a29, 'h10c26, 'h10856, 'h103bc, 'h10866, 'h10a2a, 'h10876, 'h21f8e, 'h21f8f, 'h21f8d, 'h10886, 'h10a2b, 'h10896, 'h108a6, 'h10a2c, 'h108b6, 'h108c6, 'h10a2d, 'h108d6, 'h106e6, 'h10a2e, 'h10c36, 'h106f6, 'h10706, 'h10a2f, 'h103bc, 'h10716, 'h10726, 'h10a30, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h10746, 'h10a31, 'h10756, 'h10766, 'h10a32, 'h10776, 'h10786, 'h10a33, 'h10796, 'h10c36, 'h107a6, 'h10a34, 'h107b6, 'h103bc, 'h107c6, 'h10a35, 'h107d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e6, 'h10a36, 'h107f6, 'h10806, 'h10a37, 'h10816, 'h10826, 'h10a38, 'h10836, 'h10846, 'h10a39, 'h10c36, 'h10856, 'h10866, 'h10a3a, 'h103bc, 'h10876, 'h10886, 'h10a3b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10896, 'h108a6, 'h10a3c, 'h108b6, 'h108c6, 'h10a3d, 'h108d6, 'h106e6, 'h10a3e, 'h10c46, 'h106f6, 'h10706, 'h10a3f, 'h10716, 'h103bc, 'h10726, 'h10a40, 'h10736, 'h21f8e, 'h21f8f, 'h21f8d, 'h10746, 'h10a41, 'h10756, 'h10766, 'h10a42, 'h10776, 'h10786, 'h10a43, 'h10796, 'h10c46, 'h107a6, 'h10a44, 'h107b6, 'h107c6, 'h10a45, 'h103bc, 'h107d6, 'h107e6, 'h10a46, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f6, 'h10806, 'h10a47, 'h10816, 'h10826, 'h10a48, 'h10836, 'h10846, 'h10a49, 'h10c46, 'h10856, 'h10866, 'h10a4a, 'h10876, 'h103bc, 'h10886, 'h10a4b, 'h10896, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a6, 'h10a4c, 'h108b6, 'h108c6, 'h10a4d, 'h108d6, 'h106e6, 'h10a4e, 'h10c56, 'h106f6, 'h10706, 'h10a4f, 'h10716, 'h10726, 'h10a50, 'h103bc, 'h10736, 'h10746, 'h10a51, 'h21f8e, 'h21f8f, 'h21f8d, 'h10756, 'h10766, 'h10a52, 'h10776, 'h10786, 'h10a53, 'h10796, 'h10c56, 'h107a6, 'h10a54, 'h107b6, 'h107c6, 'h10a55, 'h107d6, 'h103bc, 'h107e6, 'h10a56, 'h107f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10806, 'h10a57, 'h10816, 'h10826, 'h10a58, 'h10836, 'h10846, 'h10a59, 'h10c56, 'h10856, 'h10866, 'h10a5a, 'h10876, 'h10886, 'h10a5b, 'h103bc, 'h10896, 'h108a6, 'h10a5c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b6, 'h108c6, 'h10a5d, 'h108d6, 'h106e6, 'h10a5e, 'h10c66, 'h106f6, 'h10706, 'h10a5f, 'h10716, 'h10726, 'h10a60, 'h10736, 'h103bc, 'h10746, 'h10a61, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h10766, 'h10a62, 'h10776, 'h10786, 'h10a63, 'h10796, 'h10c66, 'h107a6, 'h10a64, 'h107b6, 'h107c6, 'h10a65, 'h107d6, 'h107e6, 'h10a66, 'h103bc, 'h107f6, 'h10806, 'h10a67, 'h21f8e, 'h21f8f, 'h21f8d, 'h10816, 'h10826, 'h10a68, 'h10836, 'h10846, 'h10a69, 'h10c66, 'h10856, 'h10866, 'h10a6a, 'h10876, 'h10886, 'h10a6b, 'h10896, 'h103bc, 'h108a6, 'h10a6c, 'h108b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c6, 'h10a6d, 'h108d6, 'h106e6, 'h10a6e, 'h10c76, 'h106f6, 'h10706, 'h10a6f, 'h10716, 'h10726, 'h10a70, 'h10736, 'h10746, 'h10a71, 'h103bc, 'h10756, 'h10766, 'h10a72, 'h21f8e, 'h21f8f, 'h21f8d, 'h10776, 'h10786, 'h10a73, 'h10796, 'h10c76, 'h107a6, 'h10a74, 'h107b6, 'h107c6, 'h10a75, 'h107d6, 'h107e6, 'h10a76, 'h107f6, 'h103bc, 'h10806, 'h10a77, 'h10816, 'h21f8e, 'h21f8f, 'h21f8d, 'h10826, 'h10a78, 'h10836, 'h10846, 'h10a79, 'h10c76, 'h10856, 'h10866, 'h10a7a, 'h10876, 'h10886, 'h10a7b, 'h10896, 'h108a6, 'h10a7c, 'h103bc, 'h108b6, 'h108c6, 'h10a7d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d6, 'h106e6, 'h10a7e, 'h10c86, 'h106f6, 'h10706, 'h10a7f, 'h10716, 'h10726, 'h10a80, 'h10736, 'h10746, 'h10a81, 'h10756, 'h103bc, 'h10766, 'h10a82, 'h10776, 'h21f8e, 'h21f8f, 'h21f8d, 'h10786, 'h10a83, 'h10796, 'h10c86, 'h107a6, 'h10a84, 'h107b6, 'h107c6, 'h10a85, 'h107d6, 'h107e6, 'h10a86, 'h107f6, 'h10806, 'h10a87, 'h103bc, 'h10816, 'h10826, 'h10a88, 'h21f8e, 'h21f8f, 'h21f8d, 'h10836, 'h10846, 'h10a89, 'h10c86, 'h10856, 'h10866, 'h10a8a, 'h10876, 'h10886, 'h10a8b, 'h10896, 'h108a6, 'h10a8c, 'h108b6, 'h103bc, 'h108c6, 'h10a8d, 'h108d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e6, 'h10a8e, 'h10c96, 'h106f6, 'h10706, 'h10a8f, 'h10716, 'h10726, 'h10a90, 'h10736, 'h10746, 'h10a91, 'h10756, 'h10766, 'h10a92, 'h103bc, 'h10776, 'h10786, 'h10a93, 'h21f8e, 'h21f8f, 'h21f8d, 'h10796, 'h10c96, 'h107a6, 'h10a94, 'h107b6, 'h107c6, 'h10a95, 'h107d6, 'h107e6, 'h10a96, 'h107f6, 'h10806, 'h10a97, 'h10816, 'h103bc, 'h10826, 'h10a98, 'h10836, 'h21f8e, 'h21f8f, 'h21f8d, 'h10846, 'h10a99, 'h10c96, 'h10856, 'h10866, 'h10a9a, 'h10876, 'h10886, 'h10a9b, 'h10896, 'h108a6, 'h10a9c, 'h108b6, 'h108c6, 'h10a9d, 'h103bc, 'h108d6, 'h106e6, 'h10a9e, 'h10ca6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f6, 'h10706, 'h10a9f, 'h10716, 'h10726, 'h10aa0, 'h10736, 'h10746, 'h10aa1, 'h10756, 'h10766, 'h10aa2, 'h10776, 'h103bc, 'h10786, 'h10aa3, 'h10796, 'h10ca6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a6, 'h10aa4, 'h107b6, 'h107c6, 'h10aa5, 'h107d6, 'h107e6, 'h10aa6, 'h107f6, 'h10806, 'h10aa7, 'h10816, 'h10826, 'h10aa8, 'h103bc, 'h10836, 'h10846, 'h10aa9, 'h10ca6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10856, 'h10866, 'h10aaa, 'h10876, 'h10886, 'h10aab, 'h10896, 'h108a6, 'h10aac, 'h108b6, 'h108c6, 'h10aad, 'h108d6, 'h103bc, 'h106e6, 'h10aae, 'h10cb6, 'h106f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h10aaf, 'h10716, 'h10726, 'h10ab0, 'h10736, 'h10746, 'h10ab1, 'h10756, 'h10766, 'h10ab2, 'h10776, 'h10786, 'h10ab3, 'h103bc, 'h10796, 'h10cb6, 'h107a6, 'h10ab4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b6, 'h107c6, 'h10ab5, 'h107d6, 'h107e6, 'h10ab6, 'h107f6, 'h10806, 'h10ab7, 'h10816, 'h10826, 'h10ab8, 'h10836, 'h103bc, 'h10846, 'h10ab9, 'h10cb6, 'h10856, 'h21f8e, 'h21f8f, 'h21f8d, 'h10866, 'h10aba, 'h10876, 'h10886, 'h10abb, 'h10896, 'h108a6, 'h10abc, 'h108b6, 'h108c6, 'h10abd, 'h108d6, 'h106e6, 'h10abe, 'h10cc6, 'h103bc, 'h106f6, 'h10706, 'h10abf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10716, 'h10726, 'h10ac0, 'h10736, 'h10746, 'h10ac1, 'h10756, 'h10766, 'h10ac2, 'h10776, 'h10786, 'h10ac3, 'h10796, 'h10cc6, 'h103bc, 'h107a6, 'h10ac4, 'h107b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c6, 'h10ac5, 'h107d6, 'h107e6, 'h10ac6, 'h107f6, 'h10806, 'h10ac7, 'h10816, 'h10826, 'h10ac8, 'h10836, 'h10846, 'h10ac9, 'h10cc6, 'h103bc, 'h10856, 'h10866, 'h10aca, 'h21f8e, 'h21f8f, 'h21f8d, 'h10876, 'h10886, 'h10acb, 'h10896, 'h108a6, 'h10acc, 'h108b6, 'h108c6, 'h10acd, 'h108d6, 'h106e6, 'h10ace, 'h10cd6, 'h106f6, 'h103bc, 'h10706, 'h10acf, 'h10716, 'h21f8e, 'h21f8f, 'h21f8d, 'h10726, 'h10ad0, 'h10736, 'h10746, 'h10ad1, 'h10756, 'h10766, 'h10ad2, 'h10776, 'h10786, 'h10ad3, 'h10796, 'h10cd6, 'h107a6, 'h10ad4, 'h103bc, 'h107b6, 'h107c6, 'h10ad5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d6, 'h107e6, 'h10ad6, 'h107f6, 'h10806, 'h10ad7, 'h10816, 'h10826, 'h10ad8, 'h10836, 'h10846, 'h10ad9, 'h10cd6, 'h10856, 'h103bc, 'h10866, 'h10ada, 'h10876, 'h21f8e, 'h21f8f, 'h21f8d, 'h10886, 'h10adb, 'h10896, 'h108a6, 'h10adc, 'h108b6, 'h108c6, 'h10add, 'h108d6, 'h106e6, 'h108de, 'h10ae6, 'h106f6, 'h10706, 'h108df, 'h103bc, 'h10716, 'h10726, 'h108e0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h10746, 'h108e1, 'h10756, 'h10766, 'h108e2, 'h10776, 'h10786, 'h108e3, 'h10796, 'h10ae6, 'h107a6, 'h108e4, 'h107b6, 'h103bc, 'h107c6, 'h108e5, 'h107d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e6, 'h108e6, 'h107f6, 'h10806, 'h108e7, 'h10816, 'h10826, 'h108e8, 'h10836, 'h10846, 'h108e9, 'h10ae6, 'h10856, 'h10866, 'h108ea, 'h103bc, 'h10876, 'h10886, 'h108eb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10896, 'h108a6, 'h108ec, 'h108b6, 'h108c6, 'h108ed, 'h108d6, 'h106e6, 'h108ee, 'h10af6, 'h106f6, 'h10706, 'h108ef, 'h10716, 'h103bc, 'h10726, 'h108f0, 'h10736, 'h21f8e, 'h21f8f, 'h21f8d, 'h10746, 'h108f1, 'h10756, 'h10766, 'h108f2, 'h10776, 'h10786, 'h108f3, 'h10796, 'h10af6, 'h107a6, 'h108f4, 'h107b6, 'h107c6, 'h108f5, 'h103bc, 'h107d6, 'h107e6, 'h108f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f6, 'h10806, 'h108f7, 'h10816, 'h10826, 'h108f8, 'h10836, 'h10846, 'h108f9, 'h10af6, 'h10856, 'h10866, 'h108fa, 'h10876, 'h103bc, 'h10886, 'h108fb, 'h10896, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a6, 'h108fc, 'h108b6, 'h108c6, 'h108fd, 'h108d6, 'h106e6, 'h108fe, 'h10b06, 'h106f6, 'h10706, 'h108ff, 'h10716, 'h10726, 'h10900, 'h103bc, 'h10736, 'h10746, 'h10901, 'h21f8e, 'h21f8f, 'h21f8d, 'h10756, 'h10766, 'h10902, 'h10776, 'h10786, 'h10903, 'h10796, 'h10b06, 'h107a6, 'h10904, 'h107b6, 'h107c6, 'h10905, 'h107d6, 'h103bc, 'h107e6, 'h10906, 'h107f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10806, 'h10907, 'h10816, 'h10826, 'h10908, 'h10836, 'h10846, 'h10909, 'h10b06, 'h10856, 'h10866, 'h1090a, 'h10876, 'h10886, 'h1090b, 'h103bc, 'h10896, 'h108a6, 'h1090c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b6, 'h108c6, 'h1090d, 'h108d6, 'h106e6, 'h1090e, 'h10b16, 'h106f6, 'h10706, 'h1090f, 'h10716, 'h10726, 'h10910, 'h10736, 'h103bc, 'h10746, 'h10911, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h10766, 'h10912, 'h10776, 'h10786, 'h10913, 'h10796, 'h10b16, 'h107a6, 'h10914, 'h107b6, 'h107c6, 'h10915, 'h107d6, 'h107e6, 'h10916, 'h103bc, 'h107f6, 'h10806, 'h10917, 'h21f8e, 'h21f8f, 'h21f8d, 'h10816, 'h10826, 'h10918, 'h10836, 'h10846, 'h10919, 'h10b16, 'h10856, 'h10866, 'h1091a, 'h10876, 'h10886, 'h1091b, 'h10896, 'h103bc, 'h108a6, 'h1091c, 'h108b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c6, 'h1091d, 'h108d6, 'h106e6, 'h1091e, 'h10b26, 'h106f6, 'h10706, 'h1091f, 'h10716, 'h10726, 'h10920, 'h10736, 'h10746, 'h10921, 'h103bc, 'h10756, 'h10766, 'h10922, 'h21f8e, 'h21f8f, 'h21f8d, 'h10776, 'h10786, 'h10923, 'h10796, 'h10b26, 'h107a6, 'h10924, 'h107b6, 'h107c6, 'h10925, 'h107d6, 'h107e6, 'h10926, 'h107f6, 'h103bc, 'h10806, 'h10927, 'h10816, 'h21f8e, 'h21f8f, 'h21f8d, 'h10826, 'h10928, 'h10836, 'h10846, 'h10929, 'h10b26, 'h10856, 'h10866, 'h1092a, 'h10876, 'h10886, 'h1092b, 'h10896, 'h108a6, 'h1092c, 'h103bc, 'h108b6, 'h108c6, 'h1092d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d6, 'h106e6, 'h1092e, 'h10b36, 'h106f6, 'h10706, 'h1092f, 'h10716, 'h10726, 'h10930, 'h10736, 'h10746, 'h10931, 'h10756, 'h103bc, 'h10766, 'h10932, 'h10776, 'h21f8e, 'h21f8f, 'h21f8d, 'h10786, 'h10933, 'h10796, 'h10b36, 'h107a6, 'h10934, 'h107b6, 'h107c6, 'h10935, 'h107d6, 'h107e6, 'h10936, 'h107f6, 'h10806, 'h10937, 'h103bc, 'h10816, 'h10826, 'h10938, 'h21f8e, 'h21f8f, 'h21f8d, 'h10836, 'h10846, 'h10939, 'h10b36, 'h10856, 'h10866, 'h1093a, 'h10876, 'h10886, 'h1093b, 'h10896, 'h108a6, 'h1093c, 'h108b6, 'h103bc, 'h108c6, 'h1093d, 'h108d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e6, 'h1093e, 'h10b46, 'h106f6, 'h10706, 'h1093f, 'h10716, 'h10726, 'h10940, 'h10736, 'h10746, 'h10941, 'h10756, 'h10766, 'h10942, 'h103bc, 'h10776, 'h10786, 'h10943, 'h21f8e, 'h21f8f, 'h21f8d, 'h10796, 'h10b46, 'h107a6, 'h10944, 'h107b6, 'h107c6, 'h10945, 'h107d6, 'h107e6, 'h10946, 'h107f6, 'h10806, 'h10947, 'h10816, 'h103bc, 'h10826, 'h10948, 'h10836, 'h21f8e, 'h21f8f, 'h21f8d, 'h10846, 'h10949, 'h10b46, 'h10856, 'h10866, 'h1094a, 'h10876, 'h10886, 'h1094b, 'h10896, 'h108a6, 'h1094c, 'h108b6, 'h108c6, 'h1094d, 'h103bc, 'h108d6, 'h106e6, 'h1094e, 'h10b56, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f6, 'h10706, 'h1094f, 'h10716, 'h10726, 'h10950, 'h10736, 'h10746, 'h10951, 'h10756, 'h10766, 'h10952, 'h10776, 'h103bc, 'h10786, 'h10953, 'h10796, 'h10b56, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a6, 'h10954, 'h107b6, 'h107c6, 'h10955, 'h107d6, 'h107e6, 'h10956, 'h107f6, 'h10806, 'h10957, 'h10816, 'h10826, 'h10958, 'h103bc, 'h10836, 'h10846, 'h10959, 'h10b56, 'h21f8e, 'h21f8f, 'h21f8d, 'h10856, 'h10866, 'h1095a, 'h10876, 'h10886, 'h1095b, 'h10896, 'h108a6, 'h1095c, 'h108b6, 'h108c6, 'h1095d, 'h108d6, 'h103bc, 'h106e6, 'h1095e, 'h10b66, 'h106f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h1095f, 'h10716, 'h10726, 'h10960, 'h10736, 'h10746, 'h10961, 'h10756, 'h10766, 'h10962, 'h10776, 'h10786, 'h10963, 'h103bc, 'h10796, 'h10b66, 'h107a6, 'h10964, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b6, 'h107c6, 'h10965, 'h107d6, 'h107e6, 'h10966, 'h107f6, 'h10806, 'h10967, 'h10816, 'h10826, 'h10968, 'h10836, 'h103bc, 'h10846, 'h10969, 'h10b66, 'h10856, 'h21f8e, 'h21f8f, 'h21f8d, 'h10866, 'h1096a, 'h10876, 'h10886, 'h1096b, 'h10896, 'h108a6, 'h1096c, 'h108b6, 'h108c6, 'h1096d, 'h108d6, 'h106e6, 'h1096e, 'h10b76, 'h103bc, 'h106f6, 'h10706, 'h1096f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10716, 'h10726, 'h10970, 'h10736, 'h10746, 'h10971, 'h10756, 'h10766, 'h10972, 'h10776, 'h10786, 'h10973, 'h10796, 'h10b76, 'h103bc, 'h107a6, 'h10974, 'h107b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c6, 'h10975, 'h107d6, 'h107e6, 'h10976, 'h107f6, 'h10806, 'h10977, 'h10816, 'h10826, 'h10978, 'h10836, 'h10846, 'h10979, 'h10b76, 'h103bc, 'h10856, 'h10866, 'h1097a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10876, 'h10886, 'h1097b, 'h10896, 'h108a6, 'h1097c, 'h108b6, 'h108c6, 'h1097d, 'h108d6, 'h106e6, 'h1097e, 'h10b86, 'h106f6, 'h103bc, 'h10706, 'h1097f, 'h10716, 'h21f8e, 'h21f8f, 'h21f8d, 'h10726, 'h10980, 'h10736, 'h10746, 'h10981, 'h10756, 'h10766, 'h10982, 'h10776, 'h10786, 'h10983, 'h10796, 'h10b86, 'h107a6, 'h10984, 'h103bc, 'h107b6, 'h107c6, 'h10985, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d6, 'h107e6, 'h10986, 'h107f6, 'h10806, 'h10987, 'h10816, 'h10826, 'h10988, 'h10836, 'h10846, 'h10989, 'h10b86, 'h10856, 'h103bc, 'h10866, 'h1098a, 'h10876, 'h21f8e, 'h21f8f, 'h21f8d, 'h10886, 'h1098b, 'h10896, 'h108a6, 'h1098c, 'h108b6, 'h108c6, 'h1098d, 'h108d6, 'h106e6, 'h1098e, 'h10b96, 'h106f6, 'h10706, 'h1098f, 'h103bc, 'h10716, 'h10726, 'h10990, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h10746, 'h10991, 'h10756, 'h10766, 'h10992, 'h10776, 'h10786, 'h10993, 'h10796, 'h10b96, 'h107a6, 'h10994, 'h107b6, 'h103bc, 'h107c6, 'h10995, 'h107d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e6, 'h10996, 'h107f6, 'h10806, 'h10997, 'h10816, 'h10826, 'h10998, 'h10836, 'h10846, 'h10999, 'h10b96, 'h10856, 'h10866, 'h1099a, 'h103bc, 'h10876, 'h10886, 'h1099b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10896, 'h108a6, 'h1099c, 'h108b6, 'h108c6, 'h1099d, 'h108d6, 'h106e6, 'h1099e, 'h10ba6, 'h106f6, 'h10706, 'h1099f, 'h10716, 'h103bc, 'h10726, 'h109a0, 'h10736, 'h21f8e, 'h21f8f, 'h21f8d, 'h10746, 'h109a1, 'h10756, 'h10766, 'h109a2, 'h10776, 'h10786, 'h109a3, 'h10796, 'h10ba6, 'h107a6, 'h109a4, 'h107b6, 'h107c6, 'h109a5, 'h103bc, 'h107d6, 'h107e6, 'h109a6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f6, 'h10806, 'h109a7, 'h10816, 'h10826, 'h109a8, 'h10836, 'h10846, 'h109a9, 'h10ba6, 'h10856, 'h10866, 'h109aa, 'h10876, 'h103bc, 'h10886, 'h109ab, 'h10896, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a6, 'h109ac, 'h108b6, 'h108c6, 'h109ad, 'h108d6, 'h106e6, 'h109ae, 'h10bb6, 'h106f6, 'h10706, 'h109af, 'h10716, 'h10726, 'h109b0, 'h103bc, 'h10736, 'h10746, 'h109b1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10756, 'h10766, 'h109b2, 'h10776, 'h10786, 'h109b3, 'h10796, 'h10bb6, 'h107a6, 'h109b4, 'h107b6, 'h107c6, 'h109b5, 'h107d6, 'h103bc, 'h107e6, 'h109b6, 'h107f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10806, 'h109b7, 'h10816, 'h10826, 'h109b8, 'h10836, 'h10846, 'h109b9, 'h10bb6, 'h10856, 'h10866, 'h109ba, 'h10876, 'h10886, 'h109bb, 'h103bc, 'h10896, 'h108a6, 'h109bc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b6, 'h108c6, 'h109bd, 'h108d6, 'h106e6, 'h109be, 'h10bc6, 'h106f6, 'h10706, 'h109bf, 'h10716, 'h10726, 'h109c0, 'h10736, 'h103bc, 'h10746, 'h109c1, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h10766, 'h109c2, 'h10776, 'h10786, 'h109c3, 'h10796, 'h10bc6, 'h107a6, 'h109c4, 'h107b6, 'h107c6, 'h109c5, 'h107d6, 'h107e6, 'h109c6, 'h103bc, 'h107f6, 'h10806, 'h109c7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10816, 'h10826, 'h109c8, 'h10836, 'h10846, 'h109c9, 'h10bc6, 'h10856, 'h10866, 'h109ca, 'h10876, 'h10886, 'h109cb, 'h10896, 'h103bc, 'h108a6, 'h109cc, 'h108b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c6, 'h109cd, 'h108d6, 'h106e6, 'h109ce, 'h10bd6, 'h106f6, 'h10706, 'h109cf, 'h10716, 'h10726, 'h109d0, 'h10736, 'h10746, 'h109d1, 'h103bc, 'h10756, 'h10766, 'h109d2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10776, 'h10786, 'h109d3, 'h10796, 'h10bd6, 'h107a6, 'h109d4, 'h107b6, 'h107c6, 'h109d5, 'h107d6, 'h107e6, 'h109d6, 'h107f6, 'h103bc, 'h10806, 'h109d7, 'h10816, 'h21f8e, 'h21f8f, 'h21f8d, 'h10826, 'h109d8, 'h10836, 'h10846, 'h109d9, 'h10bd6, 'h10856, 'h10866, 'h109da, 'h10876, 'h10886, 'h109db, 'h10896, 'h108a6, 'h109dc, 'h103bc, 'h108b6, 'h108c6, 'h109dd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d6, 'h106e6, 'h109de, 'h10be6, 'h106f6, 'h10706, 'h109df, 'h10716, 'h10726, 'h109e0, 'h10736, 'h10746, 'h109e1, 'h10756, 'h103bc, 'h10766, 'h109e2, 'h10776, 'h21f8e, 'h21f8f, 'h21f8d, 'h10786, 'h109e3, 'h10796, 'h10be6, 'h107a6, 'h109e4, 'h107b6, 'h107c6, 'h109e5, 'h107d6, 'h107e6, 'h109e6, 'h107f6, 'h10806, 'h109e7, 'h103bc, 'h10816, 'h10826, 'h109e8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10836, 'h10846, 'h109e9, 'h10be6, 'h10856, 'h10866, 'h109ea, 'h10876, 'h10886, 'h109eb, 'h10896, 'h108a6, 'h109ec, 'h108b6, 'h103bc, 'h108c6, 'h109ed, 'h108d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e6, 'h109ee, 'h10bf6, 'h106f6, 'h10706, 'h109ef, 'h10716, 'h10726, 'h109f0, 'h10736, 'h10746, 'h109f1, 'h10756, 'h10766, 'h109f2, 'h103bc, 'h10776, 'h10786, 'h109f3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10796, 'h10bf6, 'h107a6, 'h109f4, 'h107b6, 'h107c6, 'h109f5, 'h107d6, 'h107e6, 'h109f6, 'h107f6, 'h10806, 'h109f7, 'h10816, 'h103bc, 'h10826, 'h109f8, 'h10836, 'h21f8e, 'h21f8f, 'h21f8d, 'h10846, 'h109f9, 'h10bf6, 'h10856, 'h10866, 'h109fa, 'h10876, 'h10886, 'h109fb, 'h10896, 'h108a6, 'h109fc, 'h108b6, 'h108c6, 'h109fd, 'h103bc, 'h108d6, 'h106e6, 'h109fe, 'h10c06, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f6, 'h10706, 'h109ff, 'h10716, 'h10726, 'h10a00, 'h10736, 'h10746, 'h10a01, 'h10756, 'h10766, 'h10a02, 'h10776, 'h103bc, 'h10786, 'h10a03, 'h10796, 'h10c06, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a6, 'h10a04, 'h107b6, 'h107c6, 'h10a05, 'h107d6, 'h107e6, 'h10a06, 'h107f6, 'h10806, 'h10a07, 'h10816, 'h10826, 'h10a08, 'h103bc, 'h10836, 'h10846, 'h10a09, 'h10c06, 'h21f8e, 'h21f8f, 'h21f8d, 'h10856, 'h10866, 'h10a0a, 'h10876, 'h10886, 'h10a0b, 'h10896, 'h108a6, 'h10a0c, 'h108b6, 'h108c6, 'h10a0d, 'h108d6, 'h103bc, 'h106e6, 'h10a0e, 'h10c16, 'h106f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h10a0f, 'h10716, 'h10726, 'h10a10, 'h10736, 'h10746, 'h10a11, 'h10756, 'h10766, 'h10a12, 'h10776, 'h10786, 'h10a13, 'h103bc, 'h10796, 'h10c16, 'h107a6, 'h10a14, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b6, 'h107c6, 'h10a15, 'h107d6, 'h107e6, 'h10a16, 'h107f6, 'h10806, 'h10a17, 'h10816, 'h10826, 'h10a18, 'h10836, 'h103bc, 'h10846, 'h10a19, 'h10c16, 'h10856, 'h21f8e, 'h21f8f, 'h21f8d, 'h10866, 'h10a1a, 'h10876, 'h10886, 'h10a1b, 'h10896, 'h108a6, 'h10a1c, 'h108b6, 'h108c6, 'h10a1d, 'h108d6, 'h106e6, 'h10a1e, 'h10c26, 'h103bc, 'h106f6, 'h10706, 'h10a1f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10716, 'h10726, 'h10a20, 'h10736, 'h10746, 'h10a21, 'h10756, 'h10766, 'h10a22, 'h10776, 'h10786, 'h10a23, 'h10796, 'h10c26, 'h103bc, 'h107a6, 'h10a24, 'h107b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c6, 'h10a25, 'h107d6, 'h107e6, 'h10a26, 'h107f6, 'h10806, 'h10a27, 'h10816, 'h10826, 'h10a28, 'h10836, 'h10846, 'h10a29, 'h10c26, 'h103bc, 'h10856, 'h10866, 'h10a2a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10876, 'h10886, 'h10a2b, 'h10896, 'h108a6, 'h10a2c, 'h108b6, 'h108c6, 'h10a2d, 'h108d6, 'h106e6, 'h10a2e, 'h10c36, 'h106f6, 'h103bc, 'h10706, 'h10a2f, 'h10716, 'h21f8e, 'h21f8f, 'h21f8d, 'h10726, 'h10a30, 'h10736, 'h10746, 'h10a31, 'h10756, 'h10766, 'h10a32, 'h10776, 'h10786, 'h10a33, 'h10796, 'h10c36, 'h107a6, 'h10a34, 'h103bc, 'h107b6, 'h107c6, 'h10a35, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d6, 'h107e6, 'h10a36, 'h107f6, 'h10806, 'h10a37, 'h10816, 'h10826, 'h10a38, 'h10836, 'h10846, 'h10a39, 'h10c36, 'h10856, 'h103bc, 'h10866, 'h10a3a, 'h10876, 'h21f8e, 'h21f8f, 'h21f8d, 'h10886, 'h10a3b, 'h10896, 'h108a6, 'h10a3c, 'h108b6, 'h108c6, 'h10a3d, 'h108d6, 'h106e6, 'h10a3e, 'h10c46, 'h106f6, 'h10706, 'h10a3f, 'h103bc, 'h10716, 'h10726, 'h10a40, 'h21f8e, 'h21f8f, 'h21f8d, 'h10736, 'h10746, 'h10a41, 'h10756, 'h10766, 'h10a42, 'h10776, 'h10786, 'h10a43, 'h10796, 'h10c46, 'h107a6, 'h10a44, 'h107b6, 'h103bc, 'h107c6, 'h10a45, 'h107d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e6, 'h10a46, 'h107f6, 'h10806, 'h10a47, 'h10816, 'h10826, 'h10a48, 'h10836, 'h10846, 'h10a49, 'h10c46, 'h10856, 'h10866, 'h10a4a, 'h103bc, 'h10876, 'h10886, 'h10a4b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10896, 'h108a6, 'h10a4c, 'h108b6, 'h108c6, 'h10a4d, 'h108d6, 'h106e6, 'h10a4e, 'h10c56, 'h106f6, 'h10706, 'h10a4f, 'h10716, 'h103bc, 'h10726, 'h10a50, 'h10736, 'h21f8e, 'h21f8f, 'h21f8d, 'h10746, 'h10a51, 'h10756, 'h10766, 'h10a52, 'h10776, 'h10786, 'h10a53, 'h10796, 'h10c56, 'h107a6, 'h10a54, 'h107b6, 'h107c6, 'h10a55, 'h103bc, 'h107d6, 'h107e6, 'h10a56, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f6, 'h10806, 'h10a57, 'h10816, 'h10826, 'h10a58, 'h10836, 'h10846, 'h10a59, 'h10c56, 'h10856, 'h10866, 'h10a5a, 'h10876, 'h103bc, 'h10886, 'h10a5b, 'h10896, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a6, 'h10a5c, 'h108b6, 'h108c6, 'h10a5d, 'h108d6, 'h106e6, 'h10a5e, 'h10c66, 'h106f6, 'h10706, 'h10a5f, 'h10716, 'h10726, 'h10a60, 'h103bc, 'h10736, 'h10746, 'h10a61, 'h21f8e, 'h21f8f, 'h21f8d, 'h10756, 'h10766, 'h10a62, 'h10776, 'h10786, 'h10a63, 'h10796, 'h10c66, 'h107a6, 'h10a64, 'h107b6, 'h107c6, 'h10a65, 'h107d6, 'h103bc, 'h107e6, 'h10a66, 'h107f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10806, 'h10a67, 'h10816, 'h10826, 'h10a68, 'h10836, 'h10846, 'h10a69, 'h10c66, 'h10856, 'h10866, 'h10a6a, 'h10876, 'h10886, 'h10a6b, 'h103bc, 'h10896, 'h108a6, 'h10a6c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b6, 'h108c6, 'h10a6d, 'h108d6, 'h106e6, 'h10a6e, 'h10c76, 'h106f6, 'h10706, 'h10a6f, 'h10716, 'h10726, 'h10a70, 'h10736, 'h103bc, 'h10746, 'h10a71, 'h10756, 'h21f8e, 'h21f8f, 'h21f8d, 'h10766, 'h10a72, 'h10776, 'h10786, 'h10a73, 'h10796, 'h10c76, 'h107a6, 'h10a74, 'h107b6, 'h107c6, 'h10a75, 'h107d6, 'h107e6, 'h10a76, 'h103bc, 'h107f6, 'h10806, 'h10a77, 'h21f8e, 'h21f8f, 'h21f8d, 'h10816, 'h10826, 'h10a78, 'h10836, 'h10846, 'h10a79, 'h10c76, 'h10856, 'h10866, 'h10a7a, 'h10876, 'h10886, 'h10a7b, 'h10896, 'h103bc, 'h108a6, 'h10a7c, 'h108b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c6, 'h10a7d, 'h108d6, 'h106e6, 'h10a7e, 'h10c86, 'h106f6, 'h10706, 'h10a7f, 'h10716, 'h10726, 'h10a80, 'h10736, 'h10746, 'h10a81, 'h103bc, 'h10756, 'h10766, 'h10a82, 'h21f8e, 'h21f8f, 'h21f8d, 'h10776, 'h10786, 'h10a83, 'h10796, 'h10c86, 'h107a6, 'h10a84, 'h107b6, 'h107c6, 'h10a85, 'h107d6, 'h107e6, 'h10a86, 'h107f6, 'h103bc, 'h10806, 'h10a87, 'h10816, 'h21f8e, 'h21f8f, 'h21f8d, 'h10826, 'h10a88, 'h10836, 'h10846, 'h10a89, 'h10c86, 'h10856, 'h10866, 'h10a8a, 'h10876, 'h10886, 'h10a8b, 'h10896, 'h108a6, 'h10a8c, 'h103bc, 'h108b6, 'h108c6, 'h10a8d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d6, 'h106e6, 'h10a8e, 'h10c96, 'h106f6, 'h10706, 'h10a8f, 'h10716, 'h10726, 'h10a90, 'h10736, 'h10746, 'h10a91, 'h10756, 'h103bc, 'h10766, 'h10a92, 'h10776, 'h21f8e, 'h21f8f, 'h21f8d, 'h10786, 'h10a93, 'h10796, 'h10c96, 'h107a6, 'h10a94, 'h107b6, 'h107c6, 'h10a95, 'h107d6, 'h107e6, 'h10a96, 'h107f6, 'h10806, 'h10a97, 'h103bc, 'h10816, 'h10826, 'h10a98, 'h21f8e, 'h21f8f, 'h21f8d, 'h10836, 'h10846, 'h10a99, 'h10c96, 'h10856, 'h10866, 'h10a9a, 'h10876, 'h10886, 'h10a9b, 'h10896, 'h108a6, 'h10a9c, 'h108b6, 'h103bc, 'h108c6, 'h10a9d, 'h108d6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e6, 'h10a9e, 'h10ca6, 'h106f6, 'h10706, 'h10a9f, 'h10716, 'h10726, 'h10aa0, 'h10736, 'h10746, 'h10aa1, 'h10756, 'h10766, 'h10aa2, 'h103bc, 'h10776, 'h10786, 'h10aa3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10796, 'h10ca6, 'h107a6, 'h10aa4, 'h107b6, 'h107c6, 'h10aa5, 'h107d6, 'h107e6, 'h10aa6, 'h107f6, 'h10806, 'h10aa7, 'h10816, 'h103bc, 'h10826, 'h10aa8, 'h10836, 'h21f8e, 'h21f8f, 'h21f8d, 'h10846, 'h10aa9, 'h10ca6, 'h10856, 'h10866, 'h10aaa, 'h10876, 'h10886, 'h10aab, 'h10896, 'h108a6, 'h10aac, 'h108b6, 'h108c6, 'h10aad, 'h103bc, 'h108d6, 'h106e6, 'h10aae, 'h10cb6, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f6, 'h10706, 'h10aaf, 'h10716, 'h10726, 'h10ab0, 'h10736, 'h10746, 'h10ab1, 'h10756, 'h10766, 'h10ab2, 'h10776, 'h103bc, 'h10786, 'h10ab3, 'h10796, 'h10cb6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a6, 'h10ab4, 'h107b6, 'h107c6, 'h10ab5, 'h107d6, 'h107e6, 'h10ab6, 'h107f6, 'h10806, 'h10ab7, 'h10816, 'h10826, 'h10ab8, 'h103bc, 'h10836, 'h10846, 'h10ab9, 'h10cb6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10856, 'h10866, 'h10aba, 'h10876, 'h10886, 'h10abb, 'h10896, 'h108a6, 'h10abc, 'h108b6, 'h108c6, 'h10abd, 'h108d6, 'h103bc, 'h106e6, 'h10abe, 'h10cc6, 'h106f6, 'h21f8e, 'h21f8f, 'h21f8d, 'h10706, 'h10abf, 'h10716, 'h10726, 'h10ac0, 'h10736, 'h10746, 'h10ac1, 'h10756, 'h10766, 'h10ac2, 'h10776, 'h10786, 'h10ac3, 'h103bc, 'h10796, 'h10cc6, 'h107a6, 'h10ac4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b6, 'h107c6, 'h10ac5, 'h107d6, 'h107e6, 'h10ac6, 'h107f6, 'h10806, 'h10ac7, 'h10816, 'h10826, 'h10ac8, 'h10836, 'h103bc, 'h10846, 'h10ac9, 'h10cc6, 'h10856, 'h21f8e, 'h21f8f, 'h21f8d, 'h10866, 'h10aca, 'h10876, 'h10886, 'h10acb, 'h10896, 'h108a6, 'h10acc, 'h108b6, 'h108c6, 'h10acd, 'h108d6, 'h106e6, 'h10ace, 'h10cd6, 'h103bc, 'h106f6, 'h10706, 'h10acf, 'h21f8e, 'h21f8f, 'h21f8d, 'h10716, 'h10726, 'h10ad0, 'h10736, 'h10746, 'h10ad1, 'h10756, 'h10766, 'h10ad2, 'h10776, 'h10786, 'h10ad3, 'h10796, 'h10cd6, 'h103bc, 'h107a6, 'h10ad4, 'h107b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c6, 'h10ad5, 'h107d6, 'h107e6, 'h10ad6, 'h107f6, 'h10806, 'h10ad7, 'h10816, 'h10826, 'h10ad8, 'h10836, 'h10846, 'h10ad9, 'h10cd6, 'h103bc, 'h10856, 'h10866, 'h10ada, 'h21f8e, 'h21f8f, 'h21f8d, 'h10876, 'h10886, 'h10adb, 'h10896, 'h108a6, 'h10adc, 'h108b6, 'h108c6, 'h10add, 'h108d6, 'h106e7, 'h108de, 'h10ae7, 'h106f7, 'h103bc, 'h10707, 'h108df, 'h10717, 'h21f8e, 'h21f8f, 'h21f8d, 'h10727, 'h108e0, 'h10737, 'h10747, 'h108e1, 'h10757, 'h10767, 'h108e2, 'h10777, 'h10787, 'h108e3, 'h10797, 'h10ae7, 'h107a7, 'h108e4, 'h103bc, 'h107b7, 'h107c7, 'h108e5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d7, 'h107e7, 'h108e6, 'h107f7, 'h10807, 'h108e7, 'h10817, 'h10827, 'h108e8, 'h10837, 'h10847, 'h108e9, 'h10ae7, 'h10857, 'h103bc, 'h10867, 'h108ea, 'h10877, 'h21f8e, 'h21f8f, 'h21f8d, 'h10887, 'h108eb, 'h10897, 'h108a7, 'h108ec, 'h108b7, 'h108c7, 'h108ed, 'h108d7, 'h106e7, 'h108ee, 'h10af7, 'h106f7, 'h10707, 'h108ef, 'h103bc, 'h10717, 'h10727, 'h108f0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h10747, 'h108f1, 'h10757, 'h10767, 'h108f2, 'h10777, 'h10787, 'h108f3, 'h10797, 'h10af7, 'h107a7, 'h108f4, 'h107b7, 'h103bc, 'h107c7, 'h108f5, 'h107d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e7, 'h108f6, 'h107f7, 'h10807, 'h108f7, 'h10817, 'h10827, 'h108f8, 'h10837, 'h10847, 'h108f9, 'h10af7, 'h10857, 'h10867, 'h108fa, 'h103bc, 'h10877, 'h10887, 'h108fb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10897, 'h108a7, 'h108fc, 'h108b7, 'h108c7, 'h108fd, 'h108d7, 'h106e7, 'h108fe, 'h10b07, 'h106f7, 'h10707, 'h108ff, 'h10717, 'h103bc, 'h10727, 'h10900, 'h10737, 'h21f8e, 'h21f8f, 'h21f8d, 'h10747, 'h10901, 'h10757, 'h10767, 'h10902, 'h10777, 'h10787, 'h10903, 'h10797, 'h10b07, 'h107a7, 'h10904, 'h107b7, 'h107c7, 'h10905, 'h103bc, 'h107d7, 'h107e7, 'h10906, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f7, 'h10807, 'h10907, 'h10817, 'h10827, 'h10908, 'h10837, 'h10847, 'h10909, 'h10b07, 'h10857, 'h10867, 'h1090a, 'h10877, 'h103bc, 'h10887, 'h1090b, 'h10897, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a7, 'h1090c, 'h108b7, 'h108c7, 'h1090d, 'h108d7, 'h106e7, 'h1090e, 'h10b17, 'h106f7, 'h10707, 'h1090f, 'h10717, 'h10727, 'h10910, 'h103bc, 'h10737, 'h10747, 'h10911, 'h21f8e, 'h21f8f, 'h21f8d, 'h10757, 'h10767, 'h10912, 'h10777, 'h10787, 'h10913, 'h10797, 'h10b17, 'h107a7, 'h10914, 'h107b7, 'h107c7, 'h10915, 'h107d7, 'h103bc, 'h107e7, 'h10916, 'h107f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10807, 'h10917, 'h10817, 'h10827, 'h10918, 'h10837, 'h10847, 'h10919, 'h10b17, 'h10857, 'h10867, 'h1091a, 'h10877, 'h10887, 'h1091b, 'h103bc, 'h10897, 'h108a7, 'h1091c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b7, 'h108c7, 'h1091d, 'h108d7, 'h106e7, 'h1091e, 'h10b27, 'h106f7, 'h10707, 'h1091f, 'h10717, 'h10727, 'h10920, 'h10737, 'h103bc, 'h10747, 'h10921, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h10767, 'h10922, 'h10777, 'h10787, 'h10923, 'h10797, 'h10b27, 'h107a7, 'h10924, 'h107b7, 'h107c7, 'h10925, 'h107d7, 'h107e7, 'h10926, 'h103bc, 'h107f7, 'h10807, 'h10927, 'h21f8e, 'h21f8f, 'h21f8d, 'h10817, 'h10827, 'h10928, 'h10837, 'h10847, 'h10929, 'h10b27, 'h10857, 'h10867, 'h1092a, 'h10877, 'h10887, 'h1092b, 'h10897, 'h103bc, 'h108a7, 'h1092c, 'h108b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c7, 'h1092d, 'h108d7, 'h106e7, 'h1092e, 'h10b37, 'h106f7, 'h10707, 'h1092f, 'h10717, 'h10727, 'h10930, 'h10737, 'h10747, 'h10931, 'h103bc, 'h10757, 'h10767, 'h10932, 'h21f8e, 'h21f8f, 'h21f8d, 'h10777, 'h10787, 'h10933, 'h10797, 'h10b37, 'h107a7, 'h10934, 'h107b7, 'h107c7, 'h10935, 'h107d7, 'h107e7, 'h10936, 'h107f7, 'h103bc, 'h10807, 'h10937, 'h10817, 'h21f8e, 'h21f8f, 'h21f8d, 'h10827, 'h10938, 'h10837, 'h10847, 'h10939, 'h10b37, 'h10857, 'h10867, 'h1093a, 'h10877, 'h10887, 'h1093b, 'h10897, 'h108a7, 'h1093c, 'h103bc, 'h108b7, 'h108c7, 'h1093d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d7, 'h106e7, 'h1093e, 'h10b47, 'h106f7, 'h10707, 'h1093f, 'h10717, 'h10727, 'h10940, 'h10737, 'h10747, 'h10941, 'h10757, 'h103bc, 'h10767, 'h10942, 'h10777, 'h21f8e, 'h21f8f, 'h21f8d, 'h10787, 'h10943, 'h10797, 'h10b47, 'h107a7, 'h10944, 'h107b7, 'h107c7, 'h10945, 'h107d7, 'h107e7, 'h10946, 'h107f7, 'h10807, 'h10947, 'h103bc, 'h10817, 'h10827, 'h10948, 'h21f8e, 'h21f8f, 'h21f8d, 'h10837, 'h10847, 'h10949, 'h10b47, 'h10857, 'h10867, 'h1094a, 'h10877, 'h10887, 'h1094b, 'h10897, 'h108a7, 'h1094c, 'h108b7, 'h103bc, 'h108c7, 'h1094d, 'h108d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e7, 'h1094e, 'h10b57, 'h106f7, 'h10707, 'h1094f, 'h10717, 'h10727, 'h10950, 'h10737, 'h10747, 'h10951, 'h10757, 'h10767, 'h10952, 'h103bc, 'h10777, 'h10787, 'h10953, 'h21f8e, 'h21f8f, 'h21f8d, 'h10797, 'h10b57, 'h107a7, 'h10954, 'h107b7, 'h107c7, 'h10955, 'h107d7, 'h107e7, 'h10956, 'h107f7, 'h10807, 'h10957, 'h10817, 'h103bc, 'h10827, 'h10958, 'h10837, 'h21f8e, 'h21f8f, 'h21f8d, 'h10847, 'h10959, 'h10b57, 'h10857, 'h10867, 'h1095a, 'h10877, 'h10887, 'h1095b, 'h10897, 'h108a7, 'h1095c, 'h108b7, 'h108c7, 'h1095d, 'h103bc, 'h108d7, 'h106e7, 'h1095e, 'h10b67, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f7, 'h10707, 'h1095f, 'h10717, 'h10727, 'h10960, 'h10737, 'h10747, 'h10961, 'h10757, 'h10767, 'h10962, 'h10777, 'h103bc, 'h10787, 'h10963, 'h10797, 'h10b67, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a7, 'h10964, 'h107b7, 'h107c7, 'h10965, 'h107d7, 'h107e7, 'h10966, 'h107f7, 'h10807, 'h10967, 'h10817, 'h10827, 'h10968, 'h103bc, 'h10837, 'h10847, 'h10969, 'h10b67, 'h21f8e, 'h21f8f, 'h21f8d, 'h10857, 'h10867, 'h1096a, 'h10877, 'h10887, 'h1096b, 'h10897, 'h108a7, 'h1096c, 'h108b7, 'h108c7, 'h1096d, 'h108d7, 'h103bc, 'h106e7, 'h1096e, 'h10b77, 'h106f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1096f, 'h10717, 'h10727, 'h10970, 'h10737, 'h10747, 'h10971, 'h10757, 'h10767, 'h10972, 'h10777, 'h10787, 'h10973, 'h103bc, 'h10797, 'h10b77, 'h107a7, 'h10974, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b7, 'h107c7, 'h10975, 'h107d7, 'h107e7, 'h10976, 'h107f7, 'h10807, 'h10977, 'h10817, 'h10827, 'h10978, 'h10837, 'h103bc, 'h10847, 'h10979, 'h10b77, 'h10857, 'h21f8e, 'h21f8f, 'h21f8d, 'h10867, 'h1097a, 'h10877, 'h10887, 'h1097b, 'h10897, 'h108a7, 'h1097c, 'h108b7, 'h108c7, 'h1097d, 'h108d7, 'h106e7, 'h1097e, 'h10b87, 'h103bc, 'h106f7, 'h10707, 'h1097f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10717, 'h10727, 'h10980, 'h10737, 'h10747, 'h10981, 'h10757, 'h10767, 'h10982, 'h10777, 'h10787, 'h10983, 'h10797, 'h10b87, 'h103bc, 'h107a7, 'h10984, 'h107b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c7, 'h10985, 'h107d7, 'h107e7, 'h10986, 'h107f7, 'h10807, 'h10987, 'h10817, 'h10827, 'h10988, 'h10837, 'h10847, 'h10989, 'h10b87, 'h103bc, 'h10857, 'h10867, 'h1098a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10877, 'h10887, 'h1098b, 'h10897, 'h108a7, 'h1098c, 'h108b7, 'h108c7, 'h1098d, 'h108d7, 'h106e7, 'h1098e, 'h10b97, 'h106f7, 'h103bc, 'h10707, 'h1098f, 'h10717, 'h21f8e, 'h21f8f, 'h21f8d, 'h10727, 'h10990, 'h10737, 'h10747, 'h10991, 'h10757, 'h10767, 'h10992, 'h10777, 'h10787, 'h10993, 'h10797, 'h10b97, 'h107a7, 'h10994, 'h103bc, 'h107b7, 'h107c7, 'h10995, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d7, 'h107e7, 'h10996, 'h107f7, 'h10807, 'h10997, 'h10817, 'h10827, 'h10998, 'h10837, 'h10847, 'h10999, 'h10b97, 'h10857, 'h103bc, 'h10867, 'h1099a, 'h10877, 'h21f8e, 'h21f8f, 'h21f8d, 'h10887, 'h1099b, 'h10897, 'h108a7, 'h1099c, 'h108b7, 'h108c7, 'h1099d, 'h108d7, 'h106e7, 'h1099e, 'h10ba7, 'h106f7, 'h10707, 'h1099f, 'h103bc, 'h10717, 'h10727, 'h109a0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h10747, 'h109a1, 'h10757, 'h10767, 'h109a2, 'h10777, 'h10787, 'h109a3, 'h10797, 'h10ba7, 'h107a7, 'h109a4, 'h107b7, 'h103bc, 'h107c7, 'h109a5, 'h107d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e7, 'h109a6, 'h107f7, 'h10807, 'h109a7, 'h10817, 'h10827, 'h109a8, 'h10837, 'h10847, 'h109a9, 'h10ba7, 'h10857, 'h10867, 'h109aa, 'h103bc, 'h10877, 'h10887, 'h109ab, 'h21f8e, 'h21f8f, 'h21f8d, 'h10897, 'h108a7, 'h109ac, 'h108b7, 'h108c7, 'h109ad, 'h108d7, 'h106e7, 'h109ae, 'h10bb7, 'h106f7, 'h10707, 'h109af, 'h10717, 'h103bc, 'h10727, 'h109b0, 'h10737, 'h21f8e, 'h21f8f, 'h21f8d, 'h10747, 'h109b1, 'h10757, 'h10767, 'h109b2, 'h10777, 'h10787, 'h109b3, 'h10797, 'h10bb7, 'h107a7, 'h109b4, 'h107b7, 'h107c7, 'h109b5, 'h103bc, 'h107d7, 'h107e7, 'h109b6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f7, 'h10807, 'h109b7, 'h10817, 'h10827, 'h109b8, 'h10837, 'h10847, 'h109b9, 'h10bb7, 'h10857, 'h10867, 'h109ba, 'h10877, 'h103bc, 'h10887, 'h109bb, 'h10897, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a7, 'h109bc, 'h108b7, 'h108c7, 'h109bd, 'h108d7, 'h106e7, 'h109be, 'h10bc7, 'h106f7, 'h10707, 'h109bf, 'h10717, 'h10727, 'h109c0, 'h103bc, 'h10737, 'h10747, 'h109c1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10757, 'h10767, 'h109c2, 'h10777, 'h10787, 'h109c3, 'h10797, 'h10bc7, 'h107a7, 'h109c4, 'h107b7, 'h107c7, 'h109c5, 'h107d7, 'h103bc, 'h107e7, 'h109c6, 'h107f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10807, 'h109c7, 'h10817, 'h10827, 'h109c8, 'h10837, 'h10847, 'h109c9, 'h10bc7, 'h10857, 'h10867, 'h109ca, 'h10877, 'h10887, 'h109cb, 'h103bc, 'h10897, 'h108a7, 'h109cc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b7, 'h108c7, 'h109cd, 'h108d7, 'h106e7, 'h109ce, 'h10bd7, 'h106f7, 'h10707, 'h109cf, 'h10717, 'h10727, 'h109d0, 'h10737, 'h103bc, 'h10747, 'h109d1, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h10767, 'h109d2, 'h10777, 'h10787, 'h109d3, 'h10797, 'h10bd7, 'h107a7, 'h109d4, 'h107b7, 'h107c7, 'h109d5, 'h107d7, 'h107e7, 'h109d6, 'h103bc, 'h107f7, 'h10807, 'h109d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10817, 'h10827, 'h109d8, 'h10837, 'h10847, 'h109d9, 'h10bd7, 'h10857, 'h10867, 'h109da, 'h10877, 'h10887, 'h109db, 'h10897, 'h103bc, 'h108a7, 'h109dc, 'h108b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c7, 'h109dd, 'h108d7, 'h106e7, 'h109de, 'h10be7, 'h106f7, 'h10707, 'h109df, 'h10717, 'h10727, 'h109e0, 'h10737, 'h10747, 'h109e1, 'h103bc, 'h10757, 'h10767, 'h109e2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10777, 'h10787, 'h109e3, 'h10797, 'h10be7, 'h107a7, 'h109e4, 'h107b7, 'h107c7, 'h109e5, 'h107d7, 'h107e7, 'h109e6, 'h107f7, 'h103bc, 'h10807, 'h109e7, 'h10817, 'h21f8e, 'h21f8f, 'h21f8d, 'h10827, 'h109e8, 'h10837, 'h10847, 'h109e9, 'h10be7, 'h10857, 'h10867, 'h109ea, 'h10877, 'h10887, 'h109eb, 'h10897, 'h108a7, 'h109ec, 'h103bc, 'h108b7, 'h108c7, 'h109ed, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d7, 'h106e7, 'h109ee, 'h10bf7, 'h106f7, 'h10707, 'h109ef, 'h10717, 'h10727, 'h109f0, 'h10737, 'h10747, 'h109f1, 'h10757, 'h103bc, 'h10767, 'h109f2, 'h10777, 'h21f8e, 'h21f8f, 'h21f8d, 'h10787, 'h109f3, 'h10797, 'h10bf7, 'h107a7, 'h109f4, 'h107b7, 'h107c7, 'h109f5, 'h107d7, 'h107e7, 'h109f6, 'h107f7, 'h10807, 'h109f7, 'h103bc, 'h10817, 'h10827, 'h109f8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10837, 'h10847, 'h109f9, 'h10bf7, 'h10857, 'h10867, 'h109fa, 'h10877, 'h10887, 'h109fb, 'h10897, 'h108a7, 'h109fc, 'h108b7, 'h103bc, 'h108c7, 'h109fd, 'h108d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e7, 'h109fe, 'h10c07, 'h106f7, 'h10707, 'h109ff, 'h10717, 'h10727, 'h10a00, 'h10737, 'h10747, 'h10a01, 'h10757, 'h10767, 'h10a02, 'h103bc, 'h10777, 'h10787, 'h10a03, 'h21f8e, 'h21f8f, 'h21f8d, 'h10797, 'h10c07, 'h107a7, 'h10a04, 'h107b7, 'h107c7, 'h10a05, 'h107d7, 'h107e7, 'h10a06, 'h107f7, 'h10807, 'h10a07, 'h10817, 'h103bc, 'h10827, 'h10a08, 'h10837, 'h21f8e, 'h21f8f, 'h21f8d, 'h10847, 'h10a09, 'h10c07, 'h10857, 'h10867, 'h10a0a, 'h10877, 'h10887, 'h10a0b, 'h10897, 'h108a7, 'h10a0c, 'h108b7, 'h108c7, 'h10a0d, 'h103bc, 'h108d7, 'h106e7, 'h10a0e, 'h10c17, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f7, 'h10707, 'h10a0f, 'h10717, 'h10727, 'h10a10, 'h10737, 'h10747, 'h10a11, 'h10757, 'h10767, 'h10a12, 'h10777, 'h103bc, 'h10787, 'h10a13, 'h10797, 'h10c17, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a7, 'h10a14, 'h107b7, 'h107c7, 'h10a15, 'h107d7, 'h107e7, 'h10a16, 'h107f7, 'h10807, 'h10a17, 'h10817, 'h10827, 'h10a18, 'h103bc, 'h10837, 'h10847, 'h10a19, 'h10c17, 'h21f8e, 'h21f8f, 'h21f8d, 'h10857, 'h10867, 'h10a1a, 'h10877, 'h10887, 'h10a1b, 'h10897, 'h108a7, 'h10a1c, 'h108b7, 'h108c7, 'h10a1d, 'h108d7, 'h103bc, 'h106e7, 'h10a1e, 'h10c27, 'h106f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h10a1f, 'h10717, 'h10727, 'h10a20, 'h10737, 'h10747, 'h10a21, 'h10757, 'h10767, 'h10a22, 'h10777, 'h10787, 'h10a23, 'h103bc, 'h10797, 'h10c27, 'h107a7, 'h10a24, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b7, 'h107c7, 'h10a25, 'h107d7, 'h107e7, 'h10a26, 'h107f7, 'h10807, 'h10a27, 'h10817, 'h10827, 'h10a28, 'h10837, 'h103bc, 'h10847, 'h10a29, 'h10c27, 'h10857, 'h21f8e, 'h21f8f, 'h21f8d, 'h10867, 'h10a2a, 'h10877, 'h10887, 'h10a2b, 'h10897, 'h108a7, 'h10a2c, 'h108b7, 'h108c7, 'h10a2d, 'h108d7, 'h106e7, 'h10a2e, 'h10c37, 'h103bc, 'h106f7, 'h10707, 'h10a2f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10717, 'h10727, 'h10a30, 'h10737, 'h10747, 'h10a31, 'h10757, 'h10767, 'h10a32, 'h10777, 'h10787, 'h10a33, 'h10797, 'h10c37, 'h103bc, 'h107a7, 'h10a34, 'h107b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c7, 'h10a35, 'h107d7, 'h107e7, 'h10a36, 'h107f7, 'h10807, 'h10a37, 'h10817, 'h10827, 'h10a38, 'h10837, 'h10847, 'h10a39, 'h10c37, 'h103bc, 'h10857, 'h10867, 'h10a3a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10877, 'h10887, 'h10a3b, 'h10897, 'h108a7, 'h10a3c, 'h108b7, 'h108c7, 'h10a3d, 'h108d7, 'h106e7, 'h10a3e, 'h10c47, 'h106f7, 'h103bc, 'h10707, 'h10a3f, 'h10717, 'h21f8e, 'h21f8f, 'h21f8d, 'h10727, 'h10a40, 'h10737, 'h10747, 'h10a41, 'h10757, 'h10767, 'h10a42, 'h10777, 'h10787, 'h10a43, 'h10797, 'h10c47, 'h107a7, 'h10a44, 'h103bc, 'h107b7, 'h107c7, 'h10a45, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d7, 'h107e7, 'h10a46, 'h107f7, 'h10807, 'h10a47, 'h10817, 'h10827, 'h10a48, 'h10837, 'h10847, 'h10a49, 'h10c47, 'h10857, 'h103bc, 'h10867, 'h10a4a, 'h10877, 'h21f8e, 'h21f8f, 'h21f8d, 'h10887, 'h10a4b, 'h10897, 'h108a7, 'h10a4c, 'h108b7, 'h108c7, 'h10a4d, 'h108d7, 'h106e7, 'h10a4e, 'h10c57, 'h106f7, 'h10707, 'h10a4f, 'h103bc, 'h10717, 'h10727, 'h10a50, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h10747, 'h10a51, 'h10757, 'h10767, 'h10a52, 'h10777, 'h10787, 'h10a53, 'h10797, 'h10c57, 'h107a7, 'h10a54, 'h107b7, 'h103bc, 'h107c7, 'h10a55, 'h107d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e7, 'h10a56, 'h107f7, 'h10807, 'h10a57, 'h10817, 'h10827, 'h10a58, 'h10837, 'h10847, 'h10a59, 'h10c57, 'h10857, 'h10867, 'h10a5a, 'h103bc, 'h10877, 'h10887, 'h10a5b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10897, 'h108a7, 'h10a5c, 'h108b7, 'h108c7, 'h10a5d, 'h108d7, 'h106e7, 'h10a5e, 'h10c67, 'h106f7, 'h10707, 'h10a5f, 'h10717, 'h103bc, 'h10727, 'h10a60, 'h10737, 'h21f8e, 'h21f8f, 'h21f8d, 'h10747, 'h10a61, 'h10757, 'h10767, 'h10a62, 'h10777, 'h10787, 'h10a63, 'h10797, 'h10c67, 'h107a7, 'h10a64, 'h107b7, 'h107c7, 'h10a65, 'h103bc, 'h107d7, 'h107e7, 'h10a66, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f7, 'h10807, 'h10a67, 'h10817, 'h10827, 'h10a68, 'h10837, 'h10847, 'h10a69, 'h10c67, 'h10857, 'h10867, 'h10a6a, 'h10877, 'h103bc, 'h10887, 'h10a6b, 'h10897, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a7, 'h10a6c, 'h108b7, 'h108c7, 'h10a6d, 'h108d7, 'h106e7, 'h10a6e, 'h10c77, 'h106f7, 'h10707, 'h10a6f, 'h10717, 'h10727, 'h10a70, 'h103bc, 'h10737, 'h10747, 'h10a71, 'h21f8e, 'h21f8f, 'h21f8d, 'h10757, 'h10767, 'h10a72, 'h10777, 'h10787, 'h10a73, 'h10797, 'h10c77, 'h107a7, 'h10a74, 'h107b7, 'h107c7, 'h10a75, 'h107d7, 'h103bc, 'h107e7, 'h10a76, 'h107f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10807, 'h10a77, 'h10817, 'h10827, 'h10a78, 'h10837, 'h10847, 'h10a79, 'h10c77, 'h10857, 'h10867, 'h10a7a, 'h10877, 'h10887, 'h10a7b, 'h103bc, 'h10897, 'h108a7, 'h10a7c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b7, 'h108c7, 'h10a7d, 'h108d7, 'h106e7, 'h10a7e, 'h10c87, 'h106f7, 'h10707, 'h10a7f, 'h10717, 'h10727, 'h10a80, 'h10737, 'h103bc, 'h10747, 'h10a81, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h10767, 'h10a82, 'h10777, 'h10787, 'h10a83, 'h10797, 'h10c87, 'h107a7, 'h10a84, 'h107b7, 'h107c7, 'h10a85, 'h107d7, 'h107e7, 'h10a86, 'h103bc, 'h107f7, 'h10807, 'h10a87, 'h21f8e, 'h21f8f, 'h21f8d, 'h10817, 'h10827, 'h10a88, 'h10837, 'h10847, 'h10a89, 'h10c87, 'h10857, 'h10867, 'h10a8a, 'h10877, 'h10887, 'h10a8b, 'h10897, 'h103bc, 'h108a7, 'h10a8c, 'h108b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c7, 'h10a8d, 'h108d7, 'h106e7, 'h10a8e, 'h10c97, 'h106f7, 'h10707, 'h10a8f, 'h10717, 'h10727, 'h10a90, 'h10737, 'h10747, 'h10a91, 'h103bc, 'h10757, 'h10767, 'h10a92, 'h21f8e, 'h21f8f, 'h21f8d, 'h10777, 'h10787, 'h10a93, 'h10797, 'h10c97, 'h107a7, 'h10a94, 'h107b7, 'h107c7, 'h10a95, 'h107d7, 'h107e7, 'h10a96, 'h107f7, 'h103bc, 'h10807, 'h10a97, 'h10817, 'h21f8e, 'h21f8f, 'h21f8d, 'h10827, 'h10a98, 'h10837, 'h10847, 'h10a99, 'h10c97, 'h10857, 'h10867, 'h10a9a, 'h10877, 'h10887, 'h10a9b, 'h10897, 'h108a7, 'h10a9c, 'h103bc, 'h108b7, 'h108c7, 'h10a9d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d7, 'h106e7, 'h10a9e, 'h10ca7, 'h106f7, 'h10707, 'h10a9f, 'h10717, 'h10727, 'h10aa0, 'h10737, 'h10747, 'h10aa1, 'h10757, 'h103bc, 'h10767, 'h10aa2, 'h10777, 'h21f8e, 'h21f8f, 'h21f8d, 'h10787, 'h10aa3, 'h10797, 'h10ca7, 'h107a7, 'h10aa4, 'h107b7, 'h107c7, 'h10aa5, 'h107d7, 'h107e7, 'h10aa6, 'h107f7, 'h10807, 'h10aa7, 'h103bc, 'h10817, 'h10827, 'h10aa8, 'h21f8e, 'h21f8f, 'h21f8d, 'h10837, 'h10847, 'h10aa9, 'h10ca7, 'h10857, 'h10867, 'h10aaa, 'h10877, 'h10887, 'h10aab, 'h10897, 'h108a7, 'h10aac, 'h108b7, 'h103bc, 'h108c7, 'h10aad, 'h108d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e7, 'h10aae, 'h10cb7, 'h106f7, 'h10707, 'h10aaf, 'h10717, 'h10727, 'h10ab0, 'h10737, 'h10747, 'h10ab1, 'h10757, 'h10767, 'h10ab2, 'h103bc, 'h10777, 'h10787, 'h10ab3, 'h21f8e, 'h21f8f, 'h21f8d, 'h10797, 'h10cb7, 'h107a7, 'h10ab4, 'h107b7, 'h107c7, 'h10ab5, 'h107d7, 'h107e7, 'h10ab6, 'h107f7, 'h10807, 'h10ab7, 'h10817, 'h103bc, 'h10827, 'h10ab8, 'h10837, 'h21f8e, 'h21f8f, 'h21f8d, 'h10847, 'h10ab9, 'h10cb7, 'h10857, 'h10867, 'h10aba, 'h10877, 'h10887, 'h10abb, 'h10897, 'h108a7, 'h10abc, 'h108b7, 'h108c7, 'h10abd, 'h103bc, 'h108d7, 'h106e7, 'h10abe, 'h10cc7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f7, 'h10707, 'h10abf, 'h10717, 'h10727, 'h10ac0, 'h10737, 'h10747, 'h10ac1, 'h10757, 'h10767, 'h10ac2, 'h10777, 'h103bc, 'h10787, 'h10ac3, 'h10797, 'h10cc7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a7, 'h10ac4, 'h107b7, 'h107c7, 'h10ac5, 'h107d7, 'h107e7, 'h10ac6, 'h107f7, 'h10807, 'h10ac7, 'h10817, 'h10827, 'h10ac8, 'h103bc, 'h10837, 'h10847, 'h10ac9, 'h10cc7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10857, 'h10867, 'h10aca, 'h10877, 'h10887, 'h10acb, 'h10897, 'h108a7, 'h10acc, 'h108b7, 'h108c7, 'h10acd, 'h108d7, 'h103bc, 'h106e7, 'h10ace, 'h10cd7, 'h106f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h10acf, 'h10717, 'h10727, 'h10ad0, 'h10737, 'h10747, 'h10ad1, 'h10757, 'h10767, 'h10ad2, 'h10777, 'h10787, 'h10ad3, 'h103bc, 'h10797, 'h10cd7, 'h107a7, 'h10ad4, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b7, 'h107c7, 'h10ad5, 'h107d7, 'h107e7, 'h10ad6, 'h107f7, 'h10807, 'h10ad7, 'h10817, 'h10827, 'h10ad8, 'h10837, 'h103bc, 'h10847, 'h10ad9, 'h10cd7, 'h10857, 'h21f8e, 'h21f8f, 'h21f8d, 'h10867, 'h10ada, 'h10877, 'h10887, 'h10adb, 'h10897, 'h108a7, 'h10adc, 'h108b7, 'h108c7, 'h10add, 'h108d7, 'h106e7, 'h108de, 'h10ae7, 'h103bc, 'h106f7, 'h10707, 'h108df, 'h21f8e, 'h21f8f, 'h21f8d, 'h10717, 'h10727, 'h108e0, 'h10737, 'h10747, 'h108e1, 'h10757, 'h10767, 'h108e2, 'h10777, 'h10787, 'h108e3, 'h10797, 'h10ae7, 'h103bc, 'h107a7, 'h108e4, 'h107b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c7, 'h108e5, 'h107d7, 'h107e7, 'h108e6, 'h107f7, 'h10807, 'h108e7, 'h10817, 'h10827, 'h108e8, 'h10837, 'h10847, 'h108e9, 'h10ae7, 'h103bc, 'h10857, 'h10867, 'h108ea, 'h21f8e, 'h21f8f, 'h21f8d, 'h10877, 'h10887, 'h108eb, 'h10897, 'h108a7, 'h108ec, 'h108b7, 'h108c7, 'h108ed, 'h108d7, 'h106e7, 'h108ee, 'h10af7, 'h106f7, 'h103bc, 'h10707, 'h108ef, 'h10717, 'h21f8e, 'h21f8f, 'h21f8d, 'h10727, 'h108f0, 'h10737, 'h10747, 'h108f1, 'h10757, 'h10767, 'h108f2, 'h10777, 'h10787, 'h108f3, 'h10797, 'h10af7, 'h107a7, 'h108f4, 'h103bc, 'h107b7, 'h107c7, 'h108f5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d7, 'h107e7, 'h108f6, 'h107f7, 'h10807, 'h108f7, 'h10817, 'h10827, 'h108f8, 'h10837, 'h10847, 'h108f9, 'h10af7, 'h10857, 'h103bc, 'h10867, 'h108fa, 'h10877, 'h21f8e, 'h21f8f, 'h21f8d, 'h10887, 'h108fb, 'h10897, 'h108a7, 'h108fc, 'h108b7, 'h108c7, 'h108fd, 'h108d7, 'h106e7, 'h108fe, 'h10b07, 'h106f7, 'h10707, 'h108ff, 'h103bc, 'h10717, 'h10727, 'h10900, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h10747, 'h10901, 'h10757, 'h10767, 'h10902, 'h10777, 'h10787, 'h10903, 'h10797, 'h10b07, 'h107a7, 'h10904, 'h107b7, 'h103bc, 'h107c7, 'h10905, 'h107d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e7, 'h10906, 'h107f7, 'h10807, 'h10907, 'h10817, 'h10827, 'h10908, 'h10837, 'h10847, 'h10909, 'h10b07, 'h10857, 'h10867, 'h1090a, 'h103bc, 'h10877, 'h10887, 'h1090b, 'h21f8e, 'h21f8f, 'h21f8d, 'h10897, 'h108a7, 'h1090c, 'h108b7, 'h108c7, 'h1090d, 'h108d7, 'h106e7, 'h1090e, 'h10b17, 'h106f7, 'h10707, 'h1090f, 'h10717, 'h103bc, 'h10727, 'h10910, 'h10737, 'h21f8e, 'h21f8f, 'h21f8d, 'h10747, 'h10911, 'h10757, 'h10767, 'h10912, 'h10777, 'h10787, 'h10913, 'h10797, 'h10b17, 'h107a7, 'h10914, 'h107b7, 'h107c7, 'h10915, 'h103bc, 'h107d7, 'h107e7, 'h10916, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f7, 'h10807, 'h10917, 'h10817, 'h10827, 'h10918, 'h10837, 'h10847, 'h10919, 'h10b17, 'h10857, 'h10867, 'h1091a, 'h10877, 'h103bc, 'h10887, 'h1091b, 'h10897, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a7, 'h1091c, 'h108b7, 'h108c7, 'h1091d, 'h108d7, 'h106e7, 'h1091e, 'h10b27, 'h106f7, 'h10707, 'h1091f, 'h10717, 'h10727, 'h10920, 'h103bc, 'h10737, 'h10747, 'h10921, 'h21f8e, 'h21f8f, 'h21f8d, 'h10757, 'h10767, 'h10922, 'h10777, 'h10787, 'h10923, 'h10797, 'h10b27, 'h107a7, 'h10924, 'h107b7, 'h107c7, 'h10925, 'h107d7, 'h103bc, 'h107e7, 'h10926, 'h107f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10807, 'h10927, 'h10817, 'h10827, 'h10928, 'h10837, 'h10847, 'h10929, 'h10b27, 'h10857, 'h10867, 'h1092a, 'h10877, 'h10887, 'h1092b, 'h103bc, 'h10897, 'h108a7, 'h1092c, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b7, 'h108c7, 'h1092d, 'h108d7, 'h106e7, 'h1092e, 'h10b37, 'h106f7, 'h10707, 'h1092f, 'h10717, 'h10727, 'h10930, 'h10737, 'h103bc, 'h10747, 'h10931, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h10767, 'h10932, 'h10777, 'h10787, 'h10933, 'h10797, 'h10b37, 'h107a7, 'h10934, 'h107b7, 'h107c7, 'h10935, 'h107d7, 'h107e7, 'h10936, 'h103bc, 'h107f7, 'h10807, 'h10937, 'h21f8e, 'h21f8f, 'h21f8d, 'h10817, 'h10827, 'h10938, 'h10837, 'h10847, 'h10939, 'h10b37, 'h10857, 'h10867, 'h1093a, 'h10877, 'h10887, 'h1093b, 'h10897, 'h103bc, 'h108a7, 'h1093c, 'h108b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c7, 'h1093d, 'h108d7, 'h106e7, 'h1093e, 'h10b47, 'h106f7, 'h10707, 'h1093f, 'h10717, 'h10727, 'h10940, 'h10737, 'h10747, 'h10941, 'h103bc, 'h10757, 'h10767, 'h10942, 'h21f8e, 'h21f8f, 'h21f8d, 'h10777, 'h10787, 'h10943, 'h10797, 'h10b47, 'h107a7, 'h10944, 'h107b7, 'h107c7, 'h10945, 'h107d7, 'h107e7, 'h10946, 'h107f7, 'h103bc, 'h10807, 'h10947, 'h10817, 'h21f8e, 'h21f8f, 'h21f8d, 'h10827, 'h10948, 'h10837, 'h10847, 'h10949, 'h10b47, 'h10857, 'h10867, 'h1094a, 'h10877, 'h10887, 'h1094b, 'h10897, 'h108a7, 'h1094c, 'h103bc, 'h108b7, 'h108c7, 'h1094d, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d7, 'h106e7, 'h1094e, 'h10b57, 'h106f7, 'h10707, 'h1094f, 'h10717, 'h10727, 'h10950, 'h10737, 'h10747, 'h10951, 'h10757, 'h103bc, 'h10767, 'h10952, 'h10777, 'h21f8e, 'h21f8f, 'h21f8d, 'h10787, 'h10953, 'h10797, 'h10b57, 'h107a7, 'h10954, 'h107b7, 'h107c7, 'h10955, 'h107d7, 'h107e7, 'h10956, 'h107f7, 'h10807, 'h10957, 'h103bc, 'h10817, 'h10827, 'h10958, 'h21f8e, 'h21f8f, 'h21f8d, 'h10837, 'h10847, 'h10959, 'h10b57, 'h10857, 'h10867, 'h1095a, 'h10877, 'h10887, 'h1095b, 'h10897, 'h108a7, 'h1095c, 'h108b7, 'h103bc, 'h108c7, 'h1095d, 'h108d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e7, 'h1095e, 'h10b67, 'h106f7, 'h10707, 'h1095f, 'h10717, 'h10727, 'h10960, 'h10737, 'h10747, 'h10961, 'h10757, 'h10767, 'h10962, 'h103bc, 'h10777, 'h10787, 'h10963, 'h21f8e, 'h21f8f, 'h21f8d, 'h10797, 'h10b67, 'h107a7, 'h10964, 'h107b7, 'h107c7, 'h10965, 'h107d7, 'h107e7, 'h10966, 'h107f7, 'h10807, 'h10967, 'h10817, 'h103bc, 'h10827, 'h10968, 'h10837, 'h21f8e, 'h21f8f, 'h21f8d, 'h10847, 'h10969, 'h10b67, 'h10857, 'h10867, 'h1096a, 'h10877, 'h10887, 'h1096b, 'h10897, 'h108a7, 'h1096c, 'h108b7, 'h108c7, 'h1096d, 'h103bc, 'h108d7, 'h106e7, 'h1096e, 'h10b77, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f7, 'h10707, 'h1096f, 'h10717, 'h10727, 'h10970, 'h10737, 'h10747, 'h10971, 'h10757, 'h10767, 'h10972, 'h10777, 'h103bc, 'h10787, 'h10973, 'h10797, 'h10b77, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a7, 'h10974, 'h107b7, 'h107c7, 'h10975, 'h107d7, 'h107e7, 'h10976, 'h107f7, 'h10807, 'h10977, 'h10817, 'h10827, 'h10978, 'h103bc, 'h10837, 'h10847, 'h10979, 'h10b77, 'h21f8e, 'h21f8f, 'h21f8d, 'h10857, 'h10867, 'h1097a, 'h10877, 'h10887, 'h1097b, 'h10897, 'h108a7, 'h1097c, 'h108b7, 'h108c7, 'h1097d, 'h108d7, 'h103bc, 'h106e7, 'h1097e, 'h10b87, 'h106f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h1097f, 'h10717, 'h10727, 'h10980, 'h10737, 'h10747, 'h10981, 'h10757, 'h10767, 'h10982, 'h10777, 'h10787, 'h10983, 'h103bc, 'h10797, 'h10b87, 'h107a7, 'h10984, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b7, 'h107c7, 'h10985, 'h107d7, 'h107e7, 'h10986, 'h107f7, 'h10807, 'h10987, 'h10817, 'h10827, 'h10988, 'h10837, 'h103bc, 'h10847, 'h10989, 'h10b87, 'h10857, 'h21f8e, 'h21f8f, 'h21f8d, 'h10867, 'h1098a, 'h10877, 'h10887, 'h1098b, 'h10897, 'h108a7, 'h1098c, 'h108b7, 'h108c7, 'h1098d, 'h108d7, 'h106e7, 'h1098e, 'h10b97, 'h103bc, 'h106f7, 'h10707, 'h1098f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10717, 'h10727, 'h10990, 'h10737, 'h10747, 'h10991, 'h10757, 'h10767, 'h10992, 'h10777, 'h10787, 'h10993, 'h10797, 'h10b97, 'h103bc, 'h107a7, 'h10994, 'h107b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c7, 'h10995, 'h107d7, 'h107e7, 'h10996, 'h107f7, 'h10807, 'h10997, 'h10817, 'h10827, 'h10998, 'h10837, 'h10847, 'h10999, 'h10b97, 'h103bc, 'h10857, 'h10867, 'h1099a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10877, 'h10887, 'h1099b, 'h10897, 'h108a7, 'h1099c, 'h108b7, 'h108c7, 'h1099d, 'h108d7, 'h106e7, 'h1099e, 'h10ba7, 'h106f7, 'h103bc, 'h10707, 'h1099f, 'h10717, 'h21f8e, 'h21f8f, 'h21f8d, 'h10727, 'h109a0, 'h10737, 'h10747, 'h109a1, 'h10757, 'h10767, 'h109a2, 'h10777, 'h10787, 'h109a3, 'h10797, 'h10ba7, 'h107a7, 'h109a4, 'h103bc, 'h107b7, 'h107c7, 'h109a5, 'h21f8e, 'h21f8f, 'h21f8d, 'h107d7, 'h107e7, 'h109a6, 'h107f7, 'h10807, 'h109a7, 'h10817, 'h10827, 'h109a8, 'h10837, 'h10847, 'h109a9, 'h10ba7, 'h10857, 'h103bc, 'h10867, 'h109aa, 'h10877, 'h21f8e, 'h21f8f, 'h21f8d, 'h10887, 'h109ab, 'h10897, 'h108a7, 'h109ac, 'h108b7, 'h108c7, 'h109ad, 'h108d7, 'h106e7, 'h109ae, 'h10bb7, 'h106f7, 'h10707, 'h109af, 'h103bc, 'h10717, 'h10727, 'h109b0, 'h21f8e, 'h21f8f, 'h21f8d, 'h10737, 'h10747, 'h109b1, 'h10757, 'h10767, 'h109b2, 'h10777, 'h10787, 'h109b3, 'h10797, 'h10bb7, 'h107a7, 'h109b4, 'h107b7, 'h103bc, 'h107c7, 'h109b5, 'h107d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107e7, 'h109b6, 'h107f7, 'h10807, 'h109b7, 'h10817, 'h10827, 'h109b8, 'h10837, 'h10847, 'h109b9, 'h10bb7, 'h10857, 'h10867, 'h109ba, 'h103bc, 'h10877, 'h10887, 'h109bb, 'h21f8e, 'h21f8f, 'h21f8d, 'h10897, 'h108a7, 'h109bc, 'h108b7, 'h108c7, 'h109bd, 'h108d7, 'h106e7, 'h109be, 'h10bc7, 'h106f7, 'h10707, 'h109bf, 'h10717, 'h103bc, 'h10727, 'h109c0, 'h10737, 'h21f8e, 'h21f8f, 'h21f8d, 'h10747, 'h109c1, 'h10757, 'h10767, 'h109c2, 'h10777, 'h10787, 'h109c3, 'h10797, 'h10bc7, 'h107a7, 'h109c4, 'h107b7, 'h107c7, 'h109c5, 'h103bc, 'h107d7, 'h107e7, 'h109c6, 'h21f8e, 'h21f8f, 'h21f8d, 'h107f7, 'h10807, 'h109c7, 'h10817, 'h10827, 'h109c8, 'h10837, 'h10847, 'h109c9, 'h10bc7, 'h10857, 'h10867, 'h109ca, 'h10877, 'h103bc, 'h10887, 'h109cb, 'h10897, 'h21f8e, 'h21f8f, 'h21f8d, 'h108a7, 'h109cc, 'h108b7, 'h108c7, 'h109cd, 'h108d7, 'h106e7, 'h109ce, 'h10bd7, 'h106f7, 'h10707, 'h109cf, 'h10717, 'h10727, 'h109d0, 'h103bc, 'h10737, 'h10747, 'h109d1, 'h21f8e, 'h21f8f, 'h21f8d, 'h10757, 'h10767, 'h109d2, 'h10777, 'h10787, 'h109d3, 'h10797, 'h10bd7, 'h107a7, 'h109d4, 'h107b7, 'h107c7, 'h109d5, 'h107d7, 'h103bc, 'h107e7, 'h109d6, 'h107f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10807, 'h109d7, 'h10817, 'h10827, 'h109d8, 'h10837, 'h10847, 'h109d9, 'h10bd7, 'h10857, 'h10867, 'h109da, 'h10877, 'h10887, 'h109db, 'h103bc, 'h10897, 'h108a7, 'h109dc, 'h21f8e, 'h21f8f, 'h21f8d, 'h108b7, 'h108c7, 'h109dd, 'h108d7, 'h106e7, 'h109de, 'h10be7, 'h106f7, 'h10707, 'h109df, 'h10717, 'h10727, 'h109e0, 'h10737, 'h103bc, 'h10747, 'h109e1, 'h10757, 'h21f8e, 'h21f8f, 'h21f8d, 'h10767, 'h109e2, 'h10777, 'h10787, 'h109e3, 'h10797, 'h10be7, 'h107a7, 'h109e4, 'h107b7, 'h107c7, 'h109e5, 'h107d7, 'h107e7, 'h109e6, 'h103bc, 'h107f7, 'h10807, 'h109e7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10817, 'h10827, 'h109e8, 'h10837, 'h10847, 'h109e9, 'h10be7, 'h10857, 'h10867, 'h109ea, 'h10877, 'h10887, 'h109eb, 'h10897, 'h103bc, 'h108a7, 'h109ec, 'h108b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h108c7, 'h109ed, 'h108d7, 'h106e7, 'h109ee, 'h10bf7, 'h106f7, 'h10707, 'h109ef, 'h10717, 'h10727, 'h109f0, 'h10737, 'h10747, 'h109f1, 'h103bc, 'h10757, 'h10767, 'h109f2, 'h21f8e, 'h21f8f, 'h21f8d, 'h10777, 'h10787, 'h109f3, 'h10797, 'h10bf7, 'h107a7, 'h109f4, 'h107b7, 'h107c7, 'h109f5, 'h107d7, 'h107e7, 'h109f6, 'h107f7, 'h103bc, 'h10807, 'h109f7, 'h10817, 'h21f8e, 'h21f8f, 'h21f8d, 'h10827, 'h109f8, 'h10837, 'h10847, 'h109f9, 'h10bf7, 'h10857, 'h10867, 'h109fa, 'h10877, 'h10887, 'h109fb, 'h10897, 'h108a7, 'h109fc, 'h103bc, 'h108b7, 'h108c7, 'h109fd, 'h21f8e, 'h21f8f, 'h21f8d, 'h108d7, 'h106e7, 'h109fe, 'h10c07, 'h106f7, 'h10707, 'h109ff, 'h10717, 'h10727, 'h10a00, 'h10737, 'h10747, 'h10a01, 'h10757, 'h103bc, 'h10767, 'h10a02, 'h10777, 'h21f8e, 'h21f8f, 'h21f8d, 'h10787, 'h10a03, 'h10797, 'h10c07, 'h107a7, 'h10a04, 'h107b7, 'h107c7, 'h10a05, 'h107d7, 'h107e7, 'h10a06, 'h107f7, 'h10807, 'h10a07, 'h103bc, 'h10817, 'h10827, 'h10a08, 'h21f8e, 'h21f8f, 'h21f8d, 'h10837, 'h10847, 'h10a09, 'h10c07, 'h10857, 'h10867, 'h10a0a, 'h10877, 'h10887, 'h10a0b, 'h10897, 'h108a7, 'h10a0c, 'h108b7, 'h103bc, 'h108c7, 'h10a0d, 'h108d7, 'h21f8e, 'h21f8f, 'h21f8d, 'h106e7, 'h10a0e, 'h10c17, 'h106f7, 'h10707, 'h10a0f, 'h10717, 'h10727, 'h10a10, 'h10737, 'h10747, 'h10a11, 'h10757, 'h10767, 'h10a12, 'h103bc, 'h10777, 'h10787, 'h10a13, 'h21f8e, 'h21f8f, 'h21f8d, 'h10797, 'h10c17, 'h107a7, 'h10a14, 'h107b7, 'h107c7, 'h10a15, 'h107d7, 'h107e7, 'h10a16, 'h107f7, 'h10807, 'h10a17, 'h10817, 'h103bc, 'h10827, 'h10a18, 'h10837, 'h21f8e, 'h21f8f, 'h21f8d, 'h10847, 'h10a19, 'h10c17, 'h10857, 'h10867, 'h10a1a, 'h10877, 'h10887, 'h10a1b, 'h10897, 'h108a7, 'h10a1c, 'h108b7, 'h108c7, 'h10a1d, 'h103bc, 'h108d7, 'h106e7, 'h10a1e, 'h10c27, 'h21f8e, 'h21f8f, 'h21f8d, 'h106f7, 'h10707, 'h10a1f, 'h10717, 'h10727, 'h10a20, 'h10737, 'h10747, 'h10a21, 'h10757, 'h10767, 'h10a22, 'h10777, 'h103bc, 'h10787, 'h10a23, 'h10797, 'h10c27, 'h21f8e, 'h21f8f, 'h21f8d, 'h107a7, 'h10a24, 'h107b7, 'h107c7, 'h10a25, 'h107d7, 'h107e7, 'h10a26, 'h107f7, 'h10807, 'h10a27, 'h10817, 'h10827, 'h10a28, 'h103bc, 'h10837, 'h10847, 'h10a29, 'h10c27, 'h21f8e, 'h21f8f, 'h21f8d, 'h10857, 'h10867, 'h10a2a, 'h10877, 'h10887, 'h10a2b, 'h10897, 'h108a7, 'h10a2c, 'h108b7, 'h108c7, 'h10a2d, 'h108d7, 'h103bc, 'h106e7, 'h10a2e, 'h10c37, 'h106f7, 'h21f8e, 'h21f8f, 'h21f8d, 'h10707, 'h10a2f, 'h10717, 'h10727, 'h10a30, 'h10737, 'h10747, 'h10a31, 'h10757, 'h10767, 'h10a32, 'h10777, 'h10787, 'h10a33, 'h103bc, 'h10797, 'h10c37, 'h107a7, 'h10a34, 'h21f8e, 'h21f8f, 'h21f8d, 'h107b7, 'h107c7, 'h10a35, 'h107d7, 'h107e7, 'h10a36, 'h107f7, 'h10807, 'h10a37, 'h10817, 'h10827, 'h10a38, 'h10837, 'h103bc, 'h10847, 'h10a39, 'h10c37, 'h10857, 'h21f8e, 'h21f8f, 'h21f8d, 'h10867, 'h10a3a, 'h10877, 'h10887, 'h10a3b, 'h10897, 'h108a7, 'h10a3c, 'h108b7, 'h108c7, 'h10a3d, 'h108d7, 'h106e7, 'h10a3e, 'h10c47, 'h103bc, 'h106f7, 'h10707, 'h10a3f, 'h21f8e, 'h21f8f, 'h21f8d, 'h10717, 'h10727, 'h10a40, 'h10737, 'h10747, 'h10a41, 'h10757, 'h10767, 'h10a42, 'h10777, 'h10787, 'h10a43, 'h10797, 'h10c47, 'h103bc, 'h107a7, 'h10a44, 'h107b7, 'h21f8e, 'h21f8f, 'h21f8d, 'h107c7, 'h10a45, 'h107d7, 'h107e7, 'h10a46, 'h107f7, 'h10807, 'h10a47, 'h10817, 'h10827, 'h10a48, 'h10837, 'h10847, 'h10a49, 'h10c47, 'h103bc, 'h10857, 'h10867, 'h10a4a, 'h21f8e, 'h21f8f, 'h21f8d, 'h10877, 'h10887, 'h10a4b, 'h10897, 'h108a7, 'h10a4c, 'h108b7, 'h108c7, 'h10a4d, 'h108d7};
	int DATA5 [5*SIZE-1:0] = {DATA4, DATA0};
	
endpackage
